module cc_dir_ext( // @[:anonymous source@2.2]
  input  [9:0]   RW0_addr, // @[:anonymous source@3.4]
  input          RW0_clk, // @[:anonymous source@4.4]
  input  [127:0] RW0_wdata, // @[:anonymous source@5.4]
  output [127:0] RW0_rdata, // @[:anonymous source@6.4]
  input          RW0_en, // @[:anonymous source@7.4]
  input          RW0_wmode, // @[:anonymous source@8.4]
  input  [7:0]   RW0_wmask // @[:anonymous source@9.4]
);
  wire [9:0] mem_0_0_RW0_addr; // @[:anonymous source@11.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@11.4]
  wire [15:0] mem_0_0_RW0_wdata; // @[:anonymous source@11.4]
  wire [15:0] mem_0_0_RW0_rdata; // @[:anonymous source@11.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@11.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@11.4]
  wire  mem_0_0_RW0_wmask; // @[:anonymous source@11.4]
  wire [9:0] mem_0_1_RW0_addr; // @[:anonymous source@12.4]
  wire  mem_0_1_RW0_clk; // @[:anonymous source@12.4]
  wire [15:0] mem_0_1_RW0_wdata; // @[:anonymous source@12.4]
  wire [15:0] mem_0_1_RW0_rdata; // @[:anonymous source@12.4]
  wire  mem_0_1_RW0_en; // @[:anonymous source@12.4]
  wire  mem_0_1_RW0_wmode; // @[:anonymous source@12.4]
  wire  mem_0_1_RW0_wmask; // @[:anonymous source@12.4]
  wire [9:0] mem_0_2_RW0_addr; // @[:anonymous source@13.4]
  wire  mem_0_2_RW0_clk; // @[:anonymous source@13.4]
  wire [15:0] mem_0_2_RW0_wdata; // @[:anonymous source@13.4]
  wire [15:0] mem_0_2_RW0_rdata; // @[:anonymous source@13.4]
  wire  mem_0_2_RW0_en; // @[:anonymous source@13.4]
  wire  mem_0_2_RW0_wmode; // @[:anonymous source@13.4]
  wire  mem_0_2_RW0_wmask; // @[:anonymous source@13.4]
  wire [9:0] mem_0_3_RW0_addr; // @[:anonymous source@14.4]
  wire  mem_0_3_RW0_clk; // @[:anonymous source@14.4]
  wire [15:0] mem_0_3_RW0_wdata; // @[:anonymous source@14.4]
  wire [15:0] mem_0_3_RW0_rdata; // @[:anonymous source@14.4]
  wire  mem_0_3_RW0_en; // @[:anonymous source@14.4]
  wire  mem_0_3_RW0_wmode; // @[:anonymous source@14.4]
  wire  mem_0_3_RW0_wmask; // @[:anonymous source@14.4]
  wire [9:0] mem_0_4_RW0_addr; // @[:anonymous source@15.4]
  wire  mem_0_4_RW0_clk; // @[:anonymous source@15.4]
  wire [15:0] mem_0_4_RW0_wdata; // @[:anonymous source@15.4]
  wire [15:0] mem_0_4_RW0_rdata; // @[:anonymous source@15.4]
  wire  mem_0_4_RW0_en; // @[:anonymous source@15.4]
  wire  mem_0_4_RW0_wmode; // @[:anonymous source@15.4]
  wire  mem_0_4_RW0_wmask; // @[:anonymous source@15.4]
  wire [9:0] mem_0_5_RW0_addr; // @[:anonymous source@16.4]
  wire  mem_0_5_RW0_clk; // @[:anonymous source@16.4]
  wire [15:0] mem_0_5_RW0_wdata; // @[:anonymous source@16.4]
  wire [15:0] mem_0_5_RW0_rdata; // @[:anonymous source@16.4]
  wire  mem_0_5_RW0_en; // @[:anonymous source@16.4]
  wire  mem_0_5_RW0_wmode; // @[:anonymous source@16.4]
  wire  mem_0_5_RW0_wmask; // @[:anonymous source@16.4]
  wire [9:0] mem_0_6_RW0_addr; // @[:anonymous source@17.4]
  wire  mem_0_6_RW0_clk; // @[:anonymous source@17.4]
  wire [15:0] mem_0_6_RW0_wdata; // @[:anonymous source@17.4]
  wire [15:0] mem_0_6_RW0_rdata; // @[:anonymous source@17.4]
  wire  mem_0_6_RW0_en; // @[:anonymous source@17.4]
  wire  mem_0_6_RW0_wmode; // @[:anonymous source@17.4]
  wire  mem_0_6_RW0_wmask; // @[:anonymous source@17.4]
  wire [9:0] mem_0_7_RW0_addr; // @[:anonymous source@18.4]
  wire  mem_0_7_RW0_clk; // @[:anonymous source@18.4]
  wire [15:0] mem_0_7_RW0_wdata; // @[:anonymous source@18.4]
  wire [15:0] mem_0_7_RW0_rdata; // @[:anonymous source@18.4]
  wire  mem_0_7_RW0_en; // @[:anonymous source@18.4]
  wire  mem_0_7_RW0_wmode; // @[:anonymous source@18.4]
  wire  mem_0_7_RW0_wmask; // @[:anonymous source@18.4]
  wire [15:0] RW0_rdata_0_0; // @[:anonymous source@21.4]
  wire [15:0] RW0_rdata_0_1; // @[:anonymous source@28.4]
  wire [15:0] RW0_rdata_0_2; // @[:anonymous source@35.4]
  wire [15:0] RW0_rdata_0_3; // @[:anonymous source@42.4]
  wire [15:0] RW0_rdata_0_4; // @[:anonymous source@49.4]
  wire [15:0] RW0_rdata_0_5; // @[:anonymous source@56.4]
  wire [15:0] RW0_rdata_0_6; // @[:anonymous source@63.4]
  wire [15:0] RW0_rdata_0_7; // @[:anonymous source@70.4]
  wire [31:0] _GEN_0; // @[:anonymous source@75.4]
  wire [47:0] _GEN_1; // @[:anonymous source@75.4]
  wire [63:0] _GEN_2; // @[:anonymous source@75.4]
  wire [79:0] _GEN_3; // @[:anonymous source@75.4]
  wire [95:0] _GEN_4; // @[:anonymous source@75.4]
  wire [111:0] _GEN_5; // @[:anonymous source@75.4]
  wire [127:0] RW0_rdata_0; // @[:anonymous source@75.4]
  wire [31:0] _GEN_6; // @[:anonymous source@76.4]
  wire [47:0] _GEN_7; // @[:anonymous source@76.4]
  wire [63:0] _GEN_8; // @[:anonymous source@76.4]
  wire [79:0] _GEN_9; // @[:anonymous source@76.4]
  wire [95:0] _GEN_10; // @[:anonymous source@76.4]
  wire [111:0] _GEN_11; // @[:anonymous source@76.4]
  split_cc_dir_ext mem_0_0 ( // @[:anonymous source@11.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_cc_dir_ext mem_0_1 ( // @[:anonymous source@12.4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_cc_dir_ext mem_0_2 ( // @[:anonymous source@13.4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_cc_dir_ext mem_0_3 ( // @[:anonymous source@14.4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  split_cc_dir_ext mem_0_4 ( // @[:anonymous source@15.4]
    .RW0_addr(mem_0_4_RW0_addr),
    .RW0_clk(mem_0_4_RW0_clk),
    .RW0_wdata(mem_0_4_RW0_wdata),
    .RW0_rdata(mem_0_4_RW0_rdata),
    .RW0_en(mem_0_4_RW0_en),
    .RW0_wmode(mem_0_4_RW0_wmode),
    .RW0_wmask(mem_0_4_RW0_wmask)
  );
  split_cc_dir_ext mem_0_5 ( // @[:anonymous source@16.4]
    .RW0_addr(mem_0_5_RW0_addr),
    .RW0_clk(mem_0_5_RW0_clk),
    .RW0_wdata(mem_0_5_RW0_wdata),
    .RW0_rdata(mem_0_5_RW0_rdata),
    .RW0_en(mem_0_5_RW0_en),
    .RW0_wmode(mem_0_5_RW0_wmode),
    .RW0_wmask(mem_0_5_RW0_wmask)
  );
  split_cc_dir_ext mem_0_6 ( // @[:anonymous source@17.4]
    .RW0_addr(mem_0_6_RW0_addr),
    .RW0_clk(mem_0_6_RW0_clk),
    .RW0_wdata(mem_0_6_RW0_wdata),
    .RW0_rdata(mem_0_6_RW0_rdata),
    .RW0_en(mem_0_6_RW0_en),
    .RW0_wmode(mem_0_6_RW0_wmode),
    .RW0_wmask(mem_0_6_RW0_wmask)
  );
  split_cc_dir_ext mem_0_7 ( // @[:anonymous source@18.4]
    .RW0_addr(mem_0_7_RW0_addr),
    .RW0_clk(mem_0_7_RW0_clk),
    .RW0_wdata(mem_0_7_RW0_wdata),
    .RW0_rdata(mem_0_7_RW0_rdata),
    .RW0_en(mem_0_7_RW0_en),
    .RW0_wmode(mem_0_7_RW0_wmode),
    .RW0_wmask(mem_0_7_RW0_wmask)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@21.4]
  assign RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[:anonymous source@28.4]
  assign RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[:anonymous source@35.4]
  assign RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[:anonymous source@42.4]
  assign RW0_rdata_0_4 = mem_0_4_RW0_rdata; // @[:anonymous source@49.4]
  assign RW0_rdata_0_5 = mem_0_5_RW0_rdata; // @[:anonymous source@56.4]
  assign RW0_rdata_0_6 = mem_0_6_RW0_rdata; // @[:anonymous source@63.4]
  assign RW0_rdata_0_7 = mem_0_7_RW0_rdata; // @[:anonymous source@70.4]
  assign _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign _GEN_2 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign _GEN_3 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign _GEN_4 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign _GEN_5 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign RW0_rdata_0 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign _GEN_6 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@76.4]
  assign _GEN_7 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@76.4]
  assign _GEN_8 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@76.4]
  assign _GEN_9 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@76.4]
  assign _GEN_10 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@76.4]
  assign _GEN_11 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@76.4]
  assign RW0_rdata = {RW0_rdata_0_7,_GEN_5}; // @[:anonymous source@76.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@20.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@19.4]
  assign mem_0_0_RW0_wdata = RW0_wdata[15:0]; // @[:anonymous source@22.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@25.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@24.4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[:anonymous source@23.4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[:anonymous source@27.4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[:anonymous source@26.4]
  assign mem_0_1_RW0_wdata = RW0_wdata[31:16]; // @[:anonymous source@29.4]
  assign mem_0_1_RW0_en = RW0_en; // @[:anonymous source@32.4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[:anonymous source@31.4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[:anonymous source@30.4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[:anonymous source@34.4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[:anonymous source@33.4]
  assign mem_0_2_RW0_wdata = RW0_wdata[47:32]; // @[:anonymous source@36.4]
  assign mem_0_2_RW0_en = RW0_en; // @[:anonymous source@39.4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[:anonymous source@38.4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[:anonymous source@37.4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[:anonymous source@41.4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[:anonymous source@40.4]
  assign mem_0_3_RW0_wdata = RW0_wdata[63:48]; // @[:anonymous source@43.4]
  assign mem_0_3_RW0_en = RW0_en; // @[:anonymous source@46.4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[:anonymous source@45.4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[:anonymous source@44.4]
  assign mem_0_4_RW0_addr = RW0_addr; // @[:anonymous source@48.4]
  assign mem_0_4_RW0_clk = RW0_clk; // @[:anonymous source@47.4]
  assign mem_0_4_RW0_wdata = RW0_wdata[79:64]; // @[:anonymous source@50.4]
  assign mem_0_4_RW0_en = RW0_en; // @[:anonymous source@53.4]
  assign mem_0_4_RW0_wmode = RW0_wmode; // @[:anonymous source@52.4]
  assign mem_0_4_RW0_wmask = RW0_wmask[4]; // @[:anonymous source@51.4]
  assign mem_0_5_RW0_addr = RW0_addr; // @[:anonymous source@55.4]
  assign mem_0_5_RW0_clk = RW0_clk; // @[:anonymous source@54.4]
  assign mem_0_5_RW0_wdata = RW0_wdata[95:80]; // @[:anonymous source@57.4]
  assign mem_0_5_RW0_en = RW0_en; // @[:anonymous source@60.4]
  assign mem_0_5_RW0_wmode = RW0_wmode; // @[:anonymous source@59.4]
  assign mem_0_5_RW0_wmask = RW0_wmask[5]; // @[:anonymous source@58.4]
  assign mem_0_6_RW0_addr = RW0_addr; // @[:anonymous source@62.4]
  assign mem_0_6_RW0_clk = RW0_clk; // @[:anonymous source@61.4]
  assign mem_0_6_RW0_wdata = RW0_wdata[111:96]; // @[:anonymous source@64.4]
  assign mem_0_6_RW0_en = RW0_en; // @[:anonymous source@67.4]
  assign mem_0_6_RW0_wmode = RW0_wmode; // @[:anonymous source@66.4]
  assign mem_0_6_RW0_wmask = RW0_wmask[6]; // @[:anonymous source@65.4]
  assign mem_0_7_RW0_addr = RW0_addr; // @[:anonymous source@69.4]
  assign mem_0_7_RW0_clk = RW0_clk; // @[:anonymous source@68.4]
  assign mem_0_7_RW0_wdata = RW0_wdata[127:112]; // @[:anonymous source@71.4]
  assign mem_0_7_RW0_en = RW0_en; // @[:anonymous source@74.4]
  assign mem_0_7_RW0_wmode = RW0_wmode; // @[:anonymous source@73.4]
  assign mem_0_7_RW0_wmask = RW0_wmask[7]; // @[:anonymous source@72.4]
endmodule
module cc_banks_0_ext( // @[:anonymous source@78.2]
  input  [12:0] RW0_addr, // @[:anonymous source@79.4]
  input         RW0_clk, // @[:anonymous source@80.4]
  input  [63:0] RW0_wdata, // @[:anonymous source@81.4]
  output [63:0] RW0_rdata, // @[:anonymous source@82.4]
  input         RW0_en, // @[:anonymous source@83.4]
  input         RW0_wmode // @[:anonymous source@84.4]
);
  wire [12:0] mem_0_0_RW0_addr; // @[:anonymous source@86.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@86.4]
  wire [63:0] mem_0_0_RW0_wdata; // @[:anonymous source@86.4]
  wire [63:0] mem_0_0_RW0_rdata; // @[:anonymous source@86.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@86.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@86.4]
  wire [63:0] RW0_rdata_0_0; // @[:anonymous source@89.4]
  wire [63:0] RW0_rdata_0; // @[:anonymous source@93.4]
  split_cc_banks_0_ext mem_0_0 ( // @[:anonymous source@86.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@89.4]
  assign RW0_rdata_0 = RW0_rdata_0_0; // @[:anonymous source@93.4]
  assign RW0_rdata = mem_0_0_RW0_rdata; // @[:anonymous source@94.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@88.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@87.4]
  assign mem_0_0_RW0_wdata = RW0_wdata; // @[:anonymous source@90.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@92.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@91.4]
endmodule
module tag_array_ext( // @[:anonymous source@96.2]
  input  [5:0]   RW0_addr, // @[:anonymous source@97.4]
  input          RW0_clk, // @[:anonymous source@98.4]
  input  [175:0] RW0_wdata, // @[:anonymous source@99.4]
  output [175:0] RW0_rdata, // @[:anonymous source@100.4]
  input          RW0_en, // @[:anonymous source@101.4]
  input          RW0_wmode, // @[:anonymous source@102.4]
  input  [7:0]   RW0_wmask // @[:anonymous source@103.4]
);
  wire [5:0] mem_0_0_RW0_addr; // @[:anonymous source@105.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@105.4]
  wire [21:0] mem_0_0_RW0_wdata; // @[:anonymous source@105.4]
  wire [21:0] mem_0_0_RW0_rdata; // @[:anonymous source@105.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@105.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@105.4]
  wire  mem_0_0_RW0_wmask; // @[:anonymous source@105.4]
  wire [5:0] mem_0_1_RW0_addr; // @[:anonymous source@106.4]
  wire  mem_0_1_RW0_clk; // @[:anonymous source@106.4]
  wire [21:0] mem_0_1_RW0_wdata; // @[:anonymous source@106.4]
  wire [21:0] mem_0_1_RW0_rdata; // @[:anonymous source@106.4]
  wire  mem_0_1_RW0_en; // @[:anonymous source@106.4]
  wire  mem_0_1_RW0_wmode; // @[:anonymous source@106.4]
  wire  mem_0_1_RW0_wmask; // @[:anonymous source@106.4]
  wire [5:0] mem_0_2_RW0_addr; // @[:anonymous source@107.4]
  wire  mem_0_2_RW0_clk; // @[:anonymous source@107.4]
  wire [21:0] mem_0_2_RW0_wdata; // @[:anonymous source@107.4]
  wire [21:0] mem_0_2_RW0_rdata; // @[:anonymous source@107.4]
  wire  mem_0_2_RW0_en; // @[:anonymous source@107.4]
  wire  mem_0_2_RW0_wmode; // @[:anonymous source@107.4]
  wire  mem_0_2_RW0_wmask; // @[:anonymous source@107.4]
  wire [5:0] mem_0_3_RW0_addr; // @[:anonymous source@108.4]
  wire  mem_0_3_RW0_clk; // @[:anonymous source@108.4]
  wire [21:0] mem_0_3_RW0_wdata; // @[:anonymous source@108.4]
  wire [21:0] mem_0_3_RW0_rdata; // @[:anonymous source@108.4]
  wire  mem_0_3_RW0_en; // @[:anonymous source@108.4]
  wire  mem_0_3_RW0_wmode; // @[:anonymous source@108.4]
  wire  mem_0_3_RW0_wmask; // @[:anonymous source@108.4]
  wire [5:0] mem_0_4_RW0_addr; // @[:anonymous source@109.4]
  wire  mem_0_4_RW0_clk; // @[:anonymous source@109.4]
  wire [21:0] mem_0_4_RW0_wdata; // @[:anonymous source@109.4]
  wire [21:0] mem_0_4_RW0_rdata; // @[:anonymous source@109.4]
  wire  mem_0_4_RW0_en; // @[:anonymous source@109.4]
  wire  mem_0_4_RW0_wmode; // @[:anonymous source@109.4]
  wire  mem_0_4_RW0_wmask; // @[:anonymous source@109.4]
  wire [5:0] mem_0_5_RW0_addr; // @[:anonymous source@110.4]
  wire  mem_0_5_RW0_clk; // @[:anonymous source@110.4]
  wire [21:0] mem_0_5_RW0_wdata; // @[:anonymous source@110.4]
  wire [21:0] mem_0_5_RW0_rdata; // @[:anonymous source@110.4]
  wire  mem_0_5_RW0_en; // @[:anonymous source@110.4]
  wire  mem_0_5_RW0_wmode; // @[:anonymous source@110.4]
  wire  mem_0_5_RW0_wmask; // @[:anonymous source@110.4]
  wire [5:0] mem_0_6_RW0_addr; // @[:anonymous source@111.4]
  wire  mem_0_6_RW0_clk; // @[:anonymous source@111.4]
  wire [21:0] mem_0_6_RW0_wdata; // @[:anonymous source@111.4]
  wire [21:0] mem_0_6_RW0_rdata; // @[:anonymous source@111.4]
  wire  mem_0_6_RW0_en; // @[:anonymous source@111.4]
  wire  mem_0_6_RW0_wmode; // @[:anonymous source@111.4]
  wire  mem_0_6_RW0_wmask; // @[:anonymous source@111.4]
  wire [5:0] mem_0_7_RW0_addr; // @[:anonymous source@112.4]
  wire  mem_0_7_RW0_clk; // @[:anonymous source@112.4]
  wire [21:0] mem_0_7_RW0_wdata; // @[:anonymous source@112.4]
  wire [21:0] mem_0_7_RW0_rdata; // @[:anonymous source@112.4]
  wire  mem_0_7_RW0_en; // @[:anonymous source@112.4]
  wire  mem_0_7_RW0_wmode; // @[:anonymous source@112.4]
  wire  mem_0_7_RW0_wmask; // @[:anonymous source@112.4]
  wire [21:0] RW0_rdata_0_0; // @[:anonymous source@115.4]
  wire [21:0] RW0_rdata_0_1; // @[:anonymous source@122.4]
  wire [21:0] RW0_rdata_0_2; // @[:anonymous source@129.4]
  wire [21:0] RW0_rdata_0_3; // @[:anonymous source@136.4]
  wire [21:0] RW0_rdata_0_4; // @[:anonymous source@143.4]
  wire [21:0] RW0_rdata_0_5; // @[:anonymous source@150.4]
  wire [21:0] RW0_rdata_0_6; // @[:anonymous source@157.4]
  wire [21:0] RW0_rdata_0_7; // @[:anonymous source@164.4]
  wire [43:0] _GEN_0; // @[:anonymous source@169.4]
  wire [65:0] _GEN_1; // @[:anonymous source@169.4]
  wire [87:0] _GEN_2; // @[:anonymous source@169.4]
  wire [109:0] _GEN_3; // @[:anonymous source@169.4]
  wire [131:0] _GEN_4; // @[:anonymous source@169.4]
  wire [153:0] _GEN_5; // @[:anonymous source@169.4]
  wire [175:0] RW0_rdata_0; // @[:anonymous source@169.4]
  wire [43:0] _GEN_6; // @[:anonymous source@170.4]
  wire [65:0] _GEN_7; // @[:anonymous source@170.4]
  wire [87:0] _GEN_8; // @[:anonymous source@170.4]
  wire [109:0] _GEN_9; // @[:anonymous source@170.4]
  wire [131:0] _GEN_10; // @[:anonymous source@170.4]
  wire [153:0] _GEN_11; // @[:anonymous source@170.4]
  split_tag_array_ext mem_0_0 ( // @[:anonymous source@105.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_tag_array_ext mem_0_1 ( // @[:anonymous source@106.4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_tag_array_ext mem_0_2 ( // @[:anonymous source@107.4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_tag_array_ext mem_0_3 ( // @[:anonymous source@108.4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  split_tag_array_ext mem_0_4 ( // @[:anonymous source@109.4]
    .RW0_addr(mem_0_4_RW0_addr),
    .RW0_clk(mem_0_4_RW0_clk),
    .RW0_wdata(mem_0_4_RW0_wdata),
    .RW0_rdata(mem_0_4_RW0_rdata),
    .RW0_en(mem_0_4_RW0_en),
    .RW0_wmode(mem_0_4_RW0_wmode),
    .RW0_wmask(mem_0_4_RW0_wmask)
  );
  split_tag_array_ext mem_0_5 ( // @[:anonymous source@110.4]
    .RW0_addr(mem_0_5_RW0_addr),
    .RW0_clk(mem_0_5_RW0_clk),
    .RW0_wdata(mem_0_5_RW0_wdata),
    .RW0_rdata(mem_0_5_RW0_rdata),
    .RW0_en(mem_0_5_RW0_en),
    .RW0_wmode(mem_0_5_RW0_wmode),
    .RW0_wmask(mem_0_5_RW0_wmask)
  );
  split_tag_array_ext mem_0_6 ( // @[:anonymous source@111.4]
    .RW0_addr(mem_0_6_RW0_addr),
    .RW0_clk(mem_0_6_RW0_clk),
    .RW0_wdata(mem_0_6_RW0_wdata),
    .RW0_rdata(mem_0_6_RW0_rdata),
    .RW0_en(mem_0_6_RW0_en),
    .RW0_wmode(mem_0_6_RW0_wmode),
    .RW0_wmask(mem_0_6_RW0_wmask)
  );
  split_tag_array_ext mem_0_7 ( // @[:anonymous source@112.4]
    .RW0_addr(mem_0_7_RW0_addr),
    .RW0_clk(mem_0_7_RW0_clk),
    .RW0_wdata(mem_0_7_RW0_wdata),
    .RW0_rdata(mem_0_7_RW0_rdata),
    .RW0_en(mem_0_7_RW0_en),
    .RW0_wmode(mem_0_7_RW0_wmode),
    .RW0_wmask(mem_0_7_RW0_wmask)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@115.4]
  assign RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[:anonymous source@122.4]
  assign RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[:anonymous source@129.4]
  assign RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[:anonymous source@136.4]
  assign RW0_rdata_0_4 = mem_0_4_RW0_rdata; // @[:anonymous source@143.4]
  assign RW0_rdata_0_5 = mem_0_5_RW0_rdata; // @[:anonymous source@150.4]
  assign RW0_rdata_0_6 = mem_0_6_RW0_rdata; // @[:anonymous source@157.4]
  assign RW0_rdata_0_7 = mem_0_7_RW0_rdata; // @[:anonymous source@164.4]
  assign _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@169.4]
  assign _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@169.4]
  assign _GEN_2 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@169.4]
  assign _GEN_3 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@169.4]
  assign _GEN_4 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@169.4]
  assign _GEN_5 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@169.4]
  assign RW0_rdata_0 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@169.4]
  assign _GEN_6 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@170.4]
  assign _GEN_7 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@170.4]
  assign _GEN_8 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@170.4]
  assign _GEN_9 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@170.4]
  assign _GEN_10 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@170.4]
  assign _GEN_11 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@170.4]
  assign RW0_rdata = {RW0_rdata_0_7,_GEN_5}; // @[:anonymous source@170.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@114.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@113.4]
  assign mem_0_0_RW0_wdata = RW0_wdata[21:0]; // @[:anonymous source@116.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@119.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@118.4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[:anonymous source@117.4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[:anonymous source@121.4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[:anonymous source@120.4]
  assign mem_0_1_RW0_wdata = RW0_wdata[43:22]; // @[:anonymous source@123.4]
  assign mem_0_1_RW0_en = RW0_en; // @[:anonymous source@126.4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[:anonymous source@125.4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[:anonymous source@124.4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[:anonymous source@128.4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[:anonymous source@127.4]
  assign mem_0_2_RW0_wdata = RW0_wdata[65:44]; // @[:anonymous source@130.4]
  assign mem_0_2_RW0_en = RW0_en; // @[:anonymous source@133.4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[:anonymous source@132.4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[:anonymous source@131.4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[:anonymous source@135.4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[:anonymous source@134.4]
  assign mem_0_3_RW0_wdata = RW0_wdata[87:66]; // @[:anonymous source@137.4]
  assign mem_0_3_RW0_en = RW0_en; // @[:anonymous source@140.4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[:anonymous source@139.4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[:anonymous source@138.4]
  assign mem_0_4_RW0_addr = RW0_addr; // @[:anonymous source@142.4]
  assign mem_0_4_RW0_clk = RW0_clk; // @[:anonymous source@141.4]
  assign mem_0_4_RW0_wdata = RW0_wdata[109:88]; // @[:anonymous source@144.4]
  assign mem_0_4_RW0_en = RW0_en; // @[:anonymous source@147.4]
  assign mem_0_4_RW0_wmode = RW0_wmode; // @[:anonymous source@146.4]
  assign mem_0_4_RW0_wmask = RW0_wmask[4]; // @[:anonymous source@145.4]
  assign mem_0_5_RW0_addr = RW0_addr; // @[:anonymous source@149.4]
  assign mem_0_5_RW0_clk = RW0_clk; // @[:anonymous source@148.4]
  assign mem_0_5_RW0_wdata = RW0_wdata[131:110]; // @[:anonymous source@151.4]
  assign mem_0_5_RW0_en = RW0_en; // @[:anonymous source@154.4]
  assign mem_0_5_RW0_wmode = RW0_wmode; // @[:anonymous source@153.4]
  assign mem_0_5_RW0_wmask = RW0_wmask[5]; // @[:anonymous source@152.4]
  assign mem_0_6_RW0_addr = RW0_addr; // @[:anonymous source@156.4]
  assign mem_0_6_RW0_clk = RW0_clk; // @[:anonymous source@155.4]
  assign mem_0_6_RW0_wdata = RW0_wdata[153:132]; // @[:anonymous source@158.4]
  assign mem_0_6_RW0_en = RW0_en; // @[:anonymous source@161.4]
  assign mem_0_6_RW0_wmode = RW0_wmode; // @[:anonymous source@160.4]
  assign mem_0_6_RW0_wmask = RW0_wmask[6]; // @[:anonymous source@159.4]
  assign mem_0_7_RW0_addr = RW0_addr; // @[:anonymous source@163.4]
  assign mem_0_7_RW0_clk = RW0_clk; // @[:anonymous source@162.4]
  assign mem_0_7_RW0_wdata = RW0_wdata[175:154]; // @[:anonymous source@165.4]
  assign mem_0_7_RW0_en = RW0_en; // @[:anonymous source@168.4]
  assign mem_0_7_RW0_wmode = RW0_wmode; // @[:anonymous source@167.4]
  assign mem_0_7_RW0_wmask = RW0_wmask[7]; // @[:anonymous source@166.4]
endmodule
module array_0_0_ext( // @[:anonymous source@172.2]
  input  [7:0]   W0_addr, // @[:anonymous source@173.4]
  input          W0_clk, // @[:anonymous source@174.4]
  input  [127:0] W0_data, // @[:anonymous source@175.4]
  input          W0_en, // @[:anonymous source@176.4]
  input  [1:0]   W0_mask, // @[:anonymous source@177.4]
  input  [7:0]   R0_addr, // @[:anonymous source@178.4]
  input          R0_clk, // @[:anonymous source@179.4]
  output [127:0] R0_data, // @[:anonymous source@180.4]
  input          R0_en // @[:anonymous source@181.4]
);
  wire [7:0] mem_0_0_W0_addr; // @[:anonymous source@183.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@183.4]
  wire [63:0] mem_0_0_W0_data; // @[:anonymous source@183.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@183.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@183.4]
  wire [7:0] mem_0_0_R0_addr; // @[:anonymous source@183.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@183.4]
  wire [63:0] mem_0_0_R0_data; // @[:anonymous source@183.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@183.4]
  wire [7:0] mem_0_1_W0_addr; // @[:anonymous source@184.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@184.4]
  wire [63:0] mem_0_1_W0_data; // @[:anonymous source@184.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@184.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@184.4]
  wire [7:0] mem_0_1_R0_addr; // @[:anonymous source@184.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@184.4]
  wire [63:0] mem_0_1_R0_data; // @[:anonymous source@184.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@184.4]
  wire [63:0] R0_data_0_0; // @[:anonymous source@197.4]
  wire [63:0] R0_data_0_1; // @[:anonymous source@201.4]
  wire [127:0] R0_data_0; // @[:anonymous source@203.4]
  split_array_0_0_ext mem_0_0 ( // @[:anonymous source@183.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_array_0_0_ext mem_0_1 ( // @[:anonymous source@184.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@197.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@201.4]
  assign R0_data_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@203.4]
  assign R0_data = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@204.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@186.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@185.4]
  assign mem_0_0_W0_data = W0_data[63:0]; // @[:anonymous source@187.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@189.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@188.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@196.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@195.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@198.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@191.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@190.4]
  assign mem_0_1_W0_data = W0_data[127:64]; // @[:anonymous source@192.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@194.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@193.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@200.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@199.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@202.4]
endmodule
module tag_array_0_ext( // @[:anonymous source@206.2]
  input  [5:0]   RW0_addr, // @[:anonymous source@207.4]
  input          RW0_clk, // @[:anonymous source@208.4]
  input  [159:0] RW0_wdata, // @[:anonymous source@209.4]
  output [159:0] RW0_rdata, // @[:anonymous source@210.4]
  input          RW0_en, // @[:anonymous source@211.4]
  input          RW0_wmode, // @[:anonymous source@212.4]
  input  [7:0]   RW0_wmask // @[:anonymous source@213.4]
);
  wire [5:0] mem_0_0_RW0_addr; // @[:anonymous source@215.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@215.4]
  wire [19:0] mem_0_0_RW0_wdata; // @[:anonymous source@215.4]
  wire [19:0] mem_0_0_RW0_rdata; // @[:anonymous source@215.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@215.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@215.4]
  wire  mem_0_0_RW0_wmask; // @[:anonymous source@215.4]
  wire [5:0] mem_0_1_RW0_addr; // @[:anonymous source@216.4]
  wire  mem_0_1_RW0_clk; // @[:anonymous source@216.4]
  wire [19:0] mem_0_1_RW0_wdata; // @[:anonymous source@216.4]
  wire [19:0] mem_0_1_RW0_rdata; // @[:anonymous source@216.4]
  wire  mem_0_1_RW0_en; // @[:anonymous source@216.4]
  wire  mem_0_1_RW0_wmode; // @[:anonymous source@216.4]
  wire  mem_0_1_RW0_wmask; // @[:anonymous source@216.4]
  wire [5:0] mem_0_2_RW0_addr; // @[:anonymous source@217.4]
  wire  mem_0_2_RW0_clk; // @[:anonymous source@217.4]
  wire [19:0] mem_0_2_RW0_wdata; // @[:anonymous source@217.4]
  wire [19:0] mem_0_2_RW0_rdata; // @[:anonymous source@217.4]
  wire  mem_0_2_RW0_en; // @[:anonymous source@217.4]
  wire  mem_0_2_RW0_wmode; // @[:anonymous source@217.4]
  wire  mem_0_2_RW0_wmask; // @[:anonymous source@217.4]
  wire [5:0] mem_0_3_RW0_addr; // @[:anonymous source@218.4]
  wire  mem_0_3_RW0_clk; // @[:anonymous source@218.4]
  wire [19:0] mem_0_3_RW0_wdata; // @[:anonymous source@218.4]
  wire [19:0] mem_0_3_RW0_rdata; // @[:anonymous source@218.4]
  wire  mem_0_3_RW0_en; // @[:anonymous source@218.4]
  wire  mem_0_3_RW0_wmode; // @[:anonymous source@218.4]
  wire  mem_0_3_RW0_wmask; // @[:anonymous source@218.4]
  wire [5:0] mem_0_4_RW0_addr; // @[:anonymous source@219.4]
  wire  mem_0_4_RW0_clk; // @[:anonymous source@219.4]
  wire [19:0] mem_0_4_RW0_wdata; // @[:anonymous source@219.4]
  wire [19:0] mem_0_4_RW0_rdata; // @[:anonymous source@219.4]
  wire  mem_0_4_RW0_en; // @[:anonymous source@219.4]
  wire  mem_0_4_RW0_wmode; // @[:anonymous source@219.4]
  wire  mem_0_4_RW0_wmask; // @[:anonymous source@219.4]
  wire [5:0] mem_0_5_RW0_addr; // @[:anonymous source@220.4]
  wire  mem_0_5_RW0_clk; // @[:anonymous source@220.4]
  wire [19:0] mem_0_5_RW0_wdata; // @[:anonymous source@220.4]
  wire [19:0] mem_0_5_RW0_rdata; // @[:anonymous source@220.4]
  wire  mem_0_5_RW0_en; // @[:anonymous source@220.4]
  wire  mem_0_5_RW0_wmode; // @[:anonymous source@220.4]
  wire  mem_0_5_RW0_wmask; // @[:anonymous source@220.4]
  wire [5:0] mem_0_6_RW0_addr; // @[:anonymous source@221.4]
  wire  mem_0_6_RW0_clk; // @[:anonymous source@221.4]
  wire [19:0] mem_0_6_RW0_wdata; // @[:anonymous source@221.4]
  wire [19:0] mem_0_6_RW0_rdata; // @[:anonymous source@221.4]
  wire  mem_0_6_RW0_en; // @[:anonymous source@221.4]
  wire  mem_0_6_RW0_wmode; // @[:anonymous source@221.4]
  wire  mem_0_6_RW0_wmask; // @[:anonymous source@221.4]
  wire [5:0] mem_0_7_RW0_addr; // @[:anonymous source@222.4]
  wire  mem_0_7_RW0_clk; // @[:anonymous source@222.4]
  wire [19:0] mem_0_7_RW0_wdata; // @[:anonymous source@222.4]
  wire [19:0] mem_0_7_RW0_rdata; // @[:anonymous source@222.4]
  wire  mem_0_7_RW0_en; // @[:anonymous source@222.4]
  wire  mem_0_7_RW0_wmode; // @[:anonymous source@222.4]
  wire  mem_0_7_RW0_wmask; // @[:anonymous source@222.4]
  wire [19:0] RW0_rdata_0_0; // @[:anonymous source@225.4]
  wire [19:0] RW0_rdata_0_1; // @[:anonymous source@232.4]
  wire [19:0] RW0_rdata_0_2; // @[:anonymous source@239.4]
  wire [19:0] RW0_rdata_0_3; // @[:anonymous source@246.4]
  wire [19:0] RW0_rdata_0_4; // @[:anonymous source@253.4]
  wire [19:0] RW0_rdata_0_5; // @[:anonymous source@260.4]
  wire [19:0] RW0_rdata_0_6; // @[:anonymous source@267.4]
  wire [19:0] RW0_rdata_0_7; // @[:anonymous source@274.4]
  wire [39:0] _GEN_0; // @[:anonymous source@279.4]
  wire [59:0] _GEN_1; // @[:anonymous source@279.4]
  wire [79:0] _GEN_2; // @[:anonymous source@279.4]
  wire [99:0] _GEN_3; // @[:anonymous source@279.4]
  wire [119:0] _GEN_4; // @[:anonymous source@279.4]
  wire [139:0] _GEN_5; // @[:anonymous source@279.4]
  wire [159:0] RW0_rdata_0; // @[:anonymous source@279.4]
  wire [39:0] _GEN_6; // @[:anonymous source@280.4]
  wire [59:0] _GEN_7; // @[:anonymous source@280.4]
  wire [79:0] _GEN_8; // @[:anonymous source@280.4]
  wire [99:0] _GEN_9; // @[:anonymous source@280.4]
  wire [119:0] _GEN_10; // @[:anonymous source@280.4]
  wire [139:0] _GEN_11; // @[:anonymous source@280.4]
  split_tag_array_0_ext mem_0_0 ( // @[:anonymous source@215.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_1 ( // @[:anonymous source@216.4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_2 ( // @[:anonymous source@217.4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_3 ( // @[:anonymous source@218.4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_4 ( // @[:anonymous source@219.4]
    .RW0_addr(mem_0_4_RW0_addr),
    .RW0_clk(mem_0_4_RW0_clk),
    .RW0_wdata(mem_0_4_RW0_wdata),
    .RW0_rdata(mem_0_4_RW0_rdata),
    .RW0_en(mem_0_4_RW0_en),
    .RW0_wmode(mem_0_4_RW0_wmode),
    .RW0_wmask(mem_0_4_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_5 ( // @[:anonymous source@220.4]
    .RW0_addr(mem_0_5_RW0_addr),
    .RW0_clk(mem_0_5_RW0_clk),
    .RW0_wdata(mem_0_5_RW0_wdata),
    .RW0_rdata(mem_0_5_RW0_rdata),
    .RW0_en(mem_0_5_RW0_en),
    .RW0_wmode(mem_0_5_RW0_wmode),
    .RW0_wmask(mem_0_5_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_6 ( // @[:anonymous source@221.4]
    .RW0_addr(mem_0_6_RW0_addr),
    .RW0_clk(mem_0_6_RW0_clk),
    .RW0_wdata(mem_0_6_RW0_wdata),
    .RW0_rdata(mem_0_6_RW0_rdata),
    .RW0_en(mem_0_6_RW0_en),
    .RW0_wmode(mem_0_6_RW0_wmode),
    .RW0_wmask(mem_0_6_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_7 ( // @[:anonymous source@222.4]
    .RW0_addr(mem_0_7_RW0_addr),
    .RW0_clk(mem_0_7_RW0_clk),
    .RW0_wdata(mem_0_7_RW0_wdata),
    .RW0_rdata(mem_0_7_RW0_rdata),
    .RW0_en(mem_0_7_RW0_en),
    .RW0_wmode(mem_0_7_RW0_wmode),
    .RW0_wmask(mem_0_7_RW0_wmask)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@225.4]
  assign RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[:anonymous source@232.4]
  assign RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[:anonymous source@239.4]
  assign RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[:anonymous source@246.4]
  assign RW0_rdata_0_4 = mem_0_4_RW0_rdata; // @[:anonymous source@253.4]
  assign RW0_rdata_0_5 = mem_0_5_RW0_rdata; // @[:anonymous source@260.4]
  assign RW0_rdata_0_6 = mem_0_6_RW0_rdata; // @[:anonymous source@267.4]
  assign RW0_rdata_0_7 = mem_0_7_RW0_rdata; // @[:anonymous source@274.4]
  assign _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@279.4]
  assign _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@279.4]
  assign _GEN_2 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@279.4]
  assign _GEN_3 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@279.4]
  assign _GEN_4 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@279.4]
  assign _GEN_5 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@279.4]
  assign RW0_rdata_0 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@279.4]
  assign _GEN_6 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@280.4]
  assign _GEN_7 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@280.4]
  assign _GEN_8 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@280.4]
  assign _GEN_9 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@280.4]
  assign _GEN_10 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@280.4]
  assign _GEN_11 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@280.4]
  assign RW0_rdata = {RW0_rdata_0_7,_GEN_5}; // @[:anonymous source@280.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@224.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@223.4]
  assign mem_0_0_RW0_wdata = RW0_wdata[19:0]; // @[:anonymous source@226.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@229.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@228.4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[:anonymous source@227.4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[:anonymous source@231.4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[:anonymous source@230.4]
  assign mem_0_1_RW0_wdata = RW0_wdata[39:20]; // @[:anonymous source@233.4]
  assign mem_0_1_RW0_en = RW0_en; // @[:anonymous source@236.4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[:anonymous source@235.4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[:anonymous source@234.4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[:anonymous source@238.4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[:anonymous source@237.4]
  assign mem_0_2_RW0_wdata = RW0_wdata[59:40]; // @[:anonymous source@240.4]
  assign mem_0_2_RW0_en = RW0_en; // @[:anonymous source@243.4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[:anonymous source@242.4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[:anonymous source@241.4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[:anonymous source@245.4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[:anonymous source@244.4]
  assign mem_0_3_RW0_wdata = RW0_wdata[79:60]; // @[:anonymous source@247.4]
  assign mem_0_3_RW0_en = RW0_en; // @[:anonymous source@250.4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[:anonymous source@249.4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[:anonymous source@248.4]
  assign mem_0_4_RW0_addr = RW0_addr; // @[:anonymous source@252.4]
  assign mem_0_4_RW0_clk = RW0_clk; // @[:anonymous source@251.4]
  assign mem_0_4_RW0_wdata = RW0_wdata[99:80]; // @[:anonymous source@254.4]
  assign mem_0_4_RW0_en = RW0_en; // @[:anonymous source@257.4]
  assign mem_0_4_RW0_wmode = RW0_wmode; // @[:anonymous source@256.4]
  assign mem_0_4_RW0_wmask = RW0_wmask[4]; // @[:anonymous source@255.4]
  assign mem_0_5_RW0_addr = RW0_addr; // @[:anonymous source@259.4]
  assign mem_0_5_RW0_clk = RW0_clk; // @[:anonymous source@258.4]
  assign mem_0_5_RW0_wdata = RW0_wdata[119:100]; // @[:anonymous source@261.4]
  assign mem_0_5_RW0_en = RW0_en; // @[:anonymous source@264.4]
  assign mem_0_5_RW0_wmode = RW0_wmode; // @[:anonymous source@263.4]
  assign mem_0_5_RW0_wmask = RW0_wmask[5]; // @[:anonymous source@262.4]
  assign mem_0_6_RW0_addr = RW0_addr; // @[:anonymous source@266.4]
  assign mem_0_6_RW0_clk = RW0_clk; // @[:anonymous source@265.4]
  assign mem_0_6_RW0_wdata = RW0_wdata[139:120]; // @[:anonymous source@268.4]
  assign mem_0_6_RW0_en = RW0_en; // @[:anonymous source@271.4]
  assign mem_0_6_RW0_wmode = RW0_wmode; // @[:anonymous source@270.4]
  assign mem_0_6_RW0_wmask = RW0_wmask[6]; // @[:anonymous source@269.4]
  assign mem_0_7_RW0_addr = RW0_addr; // @[:anonymous source@273.4]
  assign mem_0_7_RW0_clk = RW0_clk; // @[:anonymous source@272.4]
  assign mem_0_7_RW0_wdata = RW0_wdata[159:140]; // @[:anonymous source@275.4]
  assign mem_0_7_RW0_en = RW0_en; // @[:anonymous source@278.4]
  assign mem_0_7_RW0_wmode = RW0_wmode; // @[:anonymous source@277.4]
  assign mem_0_7_RW0_wmask = RW0_wmask[7]; // @[:anonymous source@276.4]
endmodule
module dataArrayB0Way_0_ext( // @[:anonymous source@282.2]
  input  [7:0]  RW0_addr, // @[:anonymous source@283.4]
  input         RW0_clk, // @[:anonymous source@284.4]
  input  [63:0] RW0_wdata, // @[:anonymous source@285.4]
  output [63:0] RW0_rdata, // @[:anonymous source@286.4]
  input         RW0_en, // @[:anonymous source@287.4]
  input         RW0_wmode // @[:anonymous source@288.4]
);
  wire [7:0] mem_0_0_RW0_addr; // @[:anonymous source@290.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@290.4]
  wire [63:0] mem_0_0_RW0_wdata; // @[:anonymous source@290.4]
  wire [63:0] mem_0_0_RW0_rdata; // @[:anonymous source@290.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@290.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@290.4]
  wire [63:0] RW0_rdata_0_0; // @[:anonymous source@293.4]
  wire [63:0] RW0_rdata_0; // @[:anonymous source@297.4]
  split_dataArrayB0Way_0_ext mem_0_0 ( // @[:anonymous source@290.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@293.4]
  assign RW0_rdata_0 = RW0_rdata_0_0; // @[:anonymous source@297.4]
  assign RW0_rdata = mem_0_0_RW0_rdata; // @[:anonymous source@298.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@292.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@291.4]
  assign mem_0_0_RW0_wdata = RW0_wdata; // @[:anonymous source@294.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@296.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@295.4]
endmodule
module hi_us_ext( // @[:anonymous source@300.2]
  input  [6:0] W0_addr, // @[:anonymous source@301.4]
  input        W0_clk, // @[:anonymous source@302.4]
  input  [3:0] W0_data, // @[:anonymous source@303.4]
  input        W0_en, // @[:anonymous source@304.4]
  input  [3:0] W0_mask, // @[:anonymous source@305.4]
  input  [6:0] R0_addr, // @[:anonymous source@306.4]
  input        R0_clk, // @[:anonymous source@307.4]
  output [3:0] R0_data, // @[:anonymous source@308.4]
  input        R0_en // @[:anonymous source@309.4]
);
  wire [6:0] mem_0_0_W0_addr; // @[:anonymous source@311.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@311.4]
  wire  mem_0_0_W0_data; // @[:anonymous source@311.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@311.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@311.4]
  wire [6:0] mem_0_0_R0_addr; // @[:anonymous source@311.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@311.4]
  wire  mem_0_0_R0_data; // @[:anonymous source@311.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@311.4]
  wire [6:0] mem_0_1_W0_addr; // @[:anonymous source@312.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@312.4]
  wire  mem_0_1_W0_data; // @[:anonymous source@312.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@312.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@312.4]
  wire [6:0] mem_0_1_R0_addr; // @[:anonymous source@312.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@312.4]
  wire  mem_0_1_R0_data; // @[:anonymous source@312.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@312.4]
  wire [6:0] mem_0_2_W0_addr; // @[:anonymous source@313.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@313.4]
  wire  mem_0_2_W0_data; // @[:anonymous source@313.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@313.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@313.4]
  wire [6:0] mem_0_2_R0_addr; // @[:anonymous source@313.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@313.4]
  wire  mem_0_2_R0_data; // @[:anonymous source@313.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@313.4]
  wire [6:0] mem_0_3_W0_addr; // @[:anonymous source@314.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@314.4]
  wire  mem_0_3_W0_data; // @[:anonymous source@314.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@314.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@314.4]
  wire [6:0] mem_0_3_R0_addr; // @[:anonymous source@314.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@314.4]
  wire  mem_0_3_R0_data; // @[:anonymous source@314.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@314.4]
  wire  R0_data_0_0; // @[:anonymous source@337.4]
  wire  R0_data_0_1; // @[:anonymous source@341.4]
  wire  R0_data_0_2; // @[:anonymous source@345.4]
  wire  R0_data_0_3; // @[:anonymous source@349.4]
  wire [1:0] _GEN_0; // @[:anonymous source@351.4]
  wire [2:0] _GEN_1; // @[:anonymous source@351.4]
  wire [3:0] R0_data_0; // @[:anonymous source@351.4]
  wire [1:0] _GEN_2; // @[:anonymous source@352.4]
  wire [2:0] _GEN_3; // @[:anonymous source@352.4]
  split_hi_us_ext mem_0_0 ( // @[:anonymous source@311.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_hi_us_ext mem_0_1 ( // @[:anonymous source@312.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_hi_us_ext mem_0_2 ( // @[:anonymous source@313.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_hi_us_ext mem_0_3 ( // @[:anonymous source@314.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@337.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@341.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@345.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@349.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@351.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@351.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@351.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@352.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@352.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@352.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@316.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@315.4]
  assign mem_0_0_W0_data = W0_data[0]; // @[:anonymous source@317.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@319.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@318.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@336.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@335.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@338.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@321.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@320.4]
  assign mem_0_1_W0_data = W0_data[1]; // @[:anonymous source@322.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@324.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@323.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@340.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@339.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@342.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@326.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@325.4]
  assign mem_0_2_W0_data = W0_data[2]; // @[:anonymous source@327.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@329.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@328.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@344.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@343.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@346.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@331.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@330.4]
  assign mem_0_3_W0_data = W0_data[3]; // @[:anonymous source@332.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@334.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@333.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@348.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@347.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@350.4]
endmodule
module table_ext( // @[:anonymous source@354.2]
  input  [6:0]  W0_addr, // @[:anonymous source@355.4]
  input         W0_clk, // @[:anonymous source@356.4]
  input  [43:0] W0_data, // @[:anonymous source@357.4]
  input         W0_en, // @[:anonymous source@358.4]
  input  [3:0]  W0_mask, // @[:anonymous source@359.4]
  input  [6:0]  R0_addr, // @[:anonymous source@360.4]
  input         R0_clk, // @[:anonymous source@361.4]
  output [43:0] R0_data, // @[:anonymous source@362.4]
  input         R0_en // @[:anonymous source@363.4]
);
  wire [6:0] mem_0_0_W0_addr; // @[:anonymous source@365.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@365.4]
  wire [10:0] mem_0_0_W0_data; // @[:anonymous source@365.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@365.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@365.4]
  wire [6:0] mem_0_0_R0_addr; // @[:anonymous source@365.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@365.4]
  wire [10:0] mem_0_0_R0_data; // @[:anonymous source@365.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@365.4]
  wire [6:0] mem_0_1_W0_addr; // @[:anonymous source@366.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@366.4]
  wire [10:0] mem_0_1_W0_data; // @[:anonymous source@366.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@366.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@366.4]
  wire [6:0] mem_0_1_R0_addr; // @[:anonymous source@366.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@366.4]
  wire [10:0] mem_0_1_R0_data; // @[:anonymous source@366.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@366.4]
  wire [6:0] mem_0_2_W0_addr; // @[:anonymous source@367.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@367.4]
  wire [10:0] mem_0_2_W0_data; // @[:anonymous source@367.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@367.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@367.4]
  wire [6:0] mem_0_2_R0_addr; // @[:anonymous source@367.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@367.4]
  wire [10:0] mem_0_2_R0_data; // @[:anonymous source@367.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@367.4]
  wire [6:0] mem_0_3_W0_addr; // @[:anonymous source@368.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@368.4]
  wire [10:0] mem_0_3_W0_data; // @[:anonymous source@368.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@368.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@368.4]
  wire [6:0] mem_0_3_R0_addr; // @[:anonymous source@368.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@368.4]
  wire [10:0] mem_0_3_R0_data; // @[:anonymous source@368.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@368.4]
  wire [10:0] R0_data_0_0; // @[:anonymous source@391.4]
  wire [10:0] R0_data_0_1; // @[:anonymous source@395.4]
  wire [10:0] R0_data_0_2; // @[:anonymous source@399.4]
  wire [10:0] R0_data_0_3; // @[:anonymous source@403.4]
  wire [21:0] _GEN_0; // @[:anonymous source@405.4]
  wire [32:0] _GEN_1; // @[:anonymous source@405.4]
  wire [43:0] R0_data_0; // @[:anonymous source@405.4]
  wire [21:0] _GEN_2; // @[:anonymous source@406.4]
  wire [32:0] _GEN_3; // @[:anonymous source@406.4]
  split_table_ext mem_0_0 ( // @[:anonymous source@365.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_table_ext mem_0_1 ( // @[:anonymous source@366.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_table_ext mem_0_2 ( // @[:anonymous source@367.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_table_ext mem_0_3 ( // @[:anonymous source@368.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@391.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@395.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@399.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@403.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@405.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@405.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@405.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@406.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@406.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@406.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@370.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@369.4]
  assign mem_0_0_W0_data = W0_data[10:0]; // @[:anonymous source@371.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@373.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@372.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@390.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@389.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@392.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@375.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@374.4]
  assign mem_0_1_W0_data = W0_data[21:11]; // @[:anonymous source@376.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@378.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@377.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@394.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@393.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@396.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@380.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@379.4]
  assign mem_0_2_W0_data = W0_data[32:22]; // @[:anonymous source@381.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@383.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@382.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@398.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@397.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@400.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@385.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@384.4]
  assign mem_0_3_W0_data = W0_data[43:33]; // @[:anonymous source@386.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@388.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@387.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@402.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@401.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@404.4]
endmodule
module hi_us_0_ext( // @[:anonymous source@408.2]
  input  [7:0] W0_addr, // @[:anonymous source@409.4]
  input        W0_clk, // @[:anonymous source@410.4]
  input  [3:0] W0_data, // @[:anonymous source@411.4]
  input        W0_en, // @[:anonymous source@412.4]
  input  [3:0] W0_mask, // @[:anonymous source@413.4]
  input  [7:0] R0_addr, // @[:anonymous source@414.4]
  input        R0_clk, // @[:anonymous source@415.4]
  output [3:0] R0_data, // @[:anonymous source@416.4]
  input        R0_en // @[:anonymous source@417.4]
);
  wire [7:0] mem_0_0_W0_addr; // @[:anonymous source@419.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@419.4]
  wire  mem_0_0_W0_data; // @[:anonymous source@419.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@419.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@419.4]
  wire [7:0] mem_0_0_R0_addr; // @[:anonymous source@419.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@419.4]
  wire  mem_0_0_R0_data; // @[:anonymous source@419.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@419.4]
  wire [7:0] mem_0_1_W0_addr; // @[:anonymous source@420.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@420.4]
  wire  mem_0_1_W0_data; // @[:anonymous source@420.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@420.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@420.4]
  wire [7:0] mem_0_1_R0_addr; // @[:anonymous source@420.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@420.4]
  wire  mem_0_1_R0_data; // @[:anonymous source@420.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@420.4]
  wire [7:0] mem_0_2_W0_addr; // @[:anonymous source@421.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@421.4]
  wire  mem_0_2_W0_data; // @[:anonymous source@421.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@421.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@421.4]
  wire [7:0] mem_0_2_R0_addr; // @[:anonymous source@421.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@421.4]
  wire  mem_0_2_R0_data; // @[:anonymous source@421.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@421.4]
  wire [7:0] mem_0_3_W0_addr; // @[:anonymous source@422.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@422.4]
  wire  mem_0_3_W0_data; // @[:anonymous source@422.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@422.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@422.4]
  wire [7:0] mem_0_3_R0_addr; // @[:anonymous source@422.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@422.4]
  wire  mem_0_3_R0_data; // @[:anonymous source@422.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@422.4]
  wire  R0_data_0_0; // @[:anonymous source@445.4]
  wire  R0_data_0_1; // @[:anonymous source@449.4]
  wire  R0_data_0_2; // @[:anonymous source@453.4]
  wire  R0_data_0_3; // @[:anonymous source@457.4]
  wire [1:0] _GEN_0; // @[:anonymous source@459.4]
  wire [2:0] _GEN_1; // @[:anonymous source@459.4]
  wire [3:0] R0_data_0; // @[:anonymous source@459.4]
  wire [1:0] _GEN_2; // @[:anonymous source@460.4]
  wire [2:0] _GEN_3; // @[:anonymous source@460.4]
  split_hi_us_0_ext mem_0_0 ( // @[:anonymous source@419.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_hi_us_0_ext mem_0_1 ( // @[:anonymous source@420.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_hi_us_0_ext mem_0_2 ( // @[:anonymous source@421.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_hi_us_0_ext mem_0_3 ( // @[:anonymous source@422.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@445.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@449.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@453.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@457.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@459.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@459.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@459.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@460.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@460.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@460.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@424.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@423.4]
  assign mem_0_0_W0_data = W0_data[0]; // @[:anonymous source@425.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@427.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@426.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@444.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@443.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@446.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@429.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@428.4]
  assign mem_0_1_W0_data = W0_data[1]; // @[:anonymous source@430.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@432.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@431.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@448.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@447.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@450.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@434.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@433.4]
  assign mem_0_2_W0_data = W0_data[2]; // @[:anonymous source@435.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@437.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@436.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@452.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@451.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@454.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@439.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@438.4]
  assign mem_0_3_W0_data = W0_data[3]; // @[:anonymous source@440.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@442.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@441.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@456.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@455.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@458.4]
endmodule
module table_0_ext( // @[:anonymous source@462.2]
  input  [7:0]  W0_addr, // @[:anonymous source@463.4]
  input         W0_clk, // @[:anonymous source@464.4]
  input  [47:0] W0_data, // @[:anonymous source@465.4]
  input         W0_en, // @[:anonymous source@466.4]
  input  [3:0]  W0_mask, // @[:anonymous source@467.4]
  input  [7:0]  R0_addr, // @[:anonymous source@468.4]
  input         R0_clk, // @[:anonymous source@469.4]
  output [47:0] R0_data, // @[:anonymous source@470.4]
  input         R0_en // @[:anonymous source@471.4]
);
  wire [7:0] mem_0_0_W0_addr; // @[:anonymous source@473.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@473.4]
  wire [11:0] mem_0_0_W0_data; // @[:anonymous source@473.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@473.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@473.4]
  wire [7:0] mem_0_0_R0_addr; // @[:anonymous source@473.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@473.4]
  wire [11:0] mem_0_0_R0_data; // @[:anonymous source@473.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@473.4]
  wire [7:0] mem_0_1_W0_addr; // @[:anonymous source@474.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@474.4]
  wire [11:0] mem_0_1_W0_data; // @[:anonymous source@474.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@474.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@474.4]
  wire [7:0] mem_0_1_R0_addr; // @[:anonymous source@474.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@474.4]
  wire [11:0] mem_0_1_R0_data; // @[:anonymous source@474.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@474.4]
  wire [7:0] mem_0_2_W0_addr; // @[:anonymous source@475.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@475.4]
  wire [11:0] mem_0_2_W0_data; // @[:anonymous source@475.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@475.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@475.4]
  wire [7:0] mem_0_2_R0_addr; // @[:anonymous source@475.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@475.4]
  wire [11:0] mem_0_2_R0_data; // @[:anonymous source@475.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@475.4]
  wire [7:0] mem_0_3_W0_addr; // @[:anonymous source@476.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@476.4]
  wire [11:0] mem_0_3_W0_data; // @[:anonymous source@476.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@476.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@476.4]
  wire [7:0] mem_0_3_R0_addr; // @[:anonymous source@476.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@476.4]
  wire [11:0] mem_0_3_R0_data; // @[:anonymous source@476.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@476.4]
  wire [11:0] R0_data_0_0; // @[:anonymous source@499.4]
  wire [11:0] R0_data_0_1; // @[:anonymous source@503.4]
  wire [11:0] R0_data_0_2; // @[:anonymous source@507.4]
  wire [11:0] R0_data_0_3; // @[:anonymous source@511.4]
  wire [23:0] _GEN_0; // @[:anonymous source@513.4]
  wire [35:0] _GEN_1; // @[:anonymous source@513.4]
  wire [47:0] R0_data_0; // @[:anonymous source@513.4]
  wire [23:0] _GEN_2; // @[:anonymous source@514.4]
  wire [35:0] _GEN_3; // @[:anonymous source@514.4]
  split_table_0_ext mem_0_0 ( // @[:anonymous source@473.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_table_0_ext mem_0_1 ( // @[:anonymous source@474.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_table_0_ext mem_0_2 ( // @[:anonymous source@475.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_table_0_ext mem_0_3 ( // @[:anonymous source@476.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@499.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@503.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@507.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@511.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@513.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@513.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@513.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@514.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@514.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@514.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@478.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@477.4]
  assign mem_0_0_W0_data = W0_data[11:0]; // @[:anonymous source@479.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@481.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@480.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@498.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@497.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@500.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@483.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@482.4]
  assign mem_0_1_W0_data = W0_data[23:12]; // @[:anonymous source@484.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@486.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@485.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@502.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@501.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@504.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@488.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@487.4]
  assign mem_0_2_W0_data = W0_data[35:24]; // @[:anonymous source@489.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@491.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@490.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@506.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@505.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@508.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@493.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@492.4]
  assign mem_0_3_W0_data = W0_data[47:36]; // @[:anonymous source@494.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@496.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@495.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@510.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@509.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@512.4]
endmodule
module table_1_ext( // @[:anonymous source@516.2]
  input  [6:0]  W0_addr, // @[:anonymous source@517.4]
  input         W0_clk, // @[:anonymous source@518.4]
  input  [51:0] W0_data, // @[:anonymous source@519.4]
  input         W0_en, // @[:anonymous source@520.4]
  input  [3:0]  W0_mask, // @[:anonymous source@521.4]
  input  [6:0]  R0_addr, // @[:anonymous source@522.4]
  input         R0_clk, // @[:anonymous source@523.4]
  output [51:0] R0_data, // @[:anonymous source@524.4]
  input         R0_en // @[:anonymous source@525.4]
);
  wire [6:0] mem_0_0_W0_addr; // @[:anonymous source@527.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@527.4]
  wire [12:0] mem_0_0_W0_data; // @[:anonymous source@527.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@527.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@527.4]
  wire [6:0] mem_0_0_R0_addr; // @[:anonymous source@527.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@527.4]
  wire [12:0] mem_0_0_R0_data; // @[:anonymous source@527.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@527.4]
  wire [6:0] mem_0_1_W0_addr; // @[:anonymous source@528.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@528.4]
  wire [12:0] mem_0_1_W0_data; // @[:anonymous source@528.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@528.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@528.4]
  wire [6:0] mem_0_1_R0_addr; // @[:anonymous source@528.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@528.4]
  wire [12:0] mem_0_1_R0_data; // @[:anonymous source@528.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@528.4]
  wire [6:0] mem_0_2_W0_addr; // @[:anonymous source@529.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@529.4]
  wire [12:0] mem_0_2_W0_data; // @[:anonymous source@529.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@529.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@529.4]
  wire [6:0] mem_0_2_R0_addr; // @[:anonymous source@529.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@529.4]
  wire [12:0] mem_0_2_R0_data; // @[:anonymous source@529.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@529.4]
  wire [6:0] mem_0_3_W0_addr; // @[:anonymous source@530.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@530.4]
  wire [12:0] mem_0_3_W0_data; // @[:anonymous source@530.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@530.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@530.4]
  wire [6:0] mem_0_3_R0_addr; // @[:anonymous source@530.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@530.4]
  wire [12:0] mem_0_3_R0_data; // @[:anonymous source@530.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@530.4]
  wire [12:0] R0_data_0_0; // @[:anonymous source@553.4]
  wire [12:0] R0_data_0_1; // @[:anonymous source@557.4]
  wire [12:0] R0_data_0_2; // @[:anonymous source@561.4]
  wire [12:0] R0_data_0_3; // @[:anonymous source@565.4]
  wire [25:0] _GEN_0; // @[:anonymous source@567.4]
  wire [38:0] _GEN_1; // @[:anonymous source@567.4]
  wire [51:0] R0_data_0; // @[:anonymous source@567.4]
  wire [25:0] _GEN_2; // @[:anonymous source@568.4]
  wire [38:0] _GEN_3; // @[:anonymous source@568.4]
  split_table_1_ext mem_0_0 ( // @[:anonymous source@527.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_table_1_ext mem_0_1 ( // @[:anonymous source@528.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_table_1_ext mem_0_2 ( // @[:anonymous source@529.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_table_1_ext mem_0_3 ( // @[:anonymous source@530.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@553.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@557.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@561.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@565.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@567.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@567.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@567.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@568.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@568.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@568.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@532.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@531.4]
  assign mem_0_0_W0_data = W0_data[12:0]; // @[:anonymous source@533.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@535.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@534.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@552.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@551.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@554.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@537.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@536.4]
  assign mem_0_1_W0_data = W0_data[25:13]; // @[:anonymous source@538.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@540.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@539.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@556.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@555.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@558.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@542.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@541.4]
  assign mem_0_2_W0_data = W0_data[38:26]; // @[:anonymous source@543.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@545.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@544.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@560.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@559.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@562.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@547.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@546.4]
  assign mem_0_3_W0_data = W0_data[51:39]; // @[:anonymous source@548.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@550.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@549.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@564.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@563.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@566.4]
endmodule
module meta_0_ext( // @[:anonymous source@570.2]
  input  [6:0]   W0_addr, // @[:anonymous source@571.4]
  input          W0_clk, // @[:anonymous source@572.4]
  input  [119:0] W0_data, // @[:anonymous source@573.4]
  input          W0_en, // @[:anonymous source@574.4]
  input  [3:0]   W0_mask, // @[:anonymous source@575.4]
  input  [6:0]   R0_addr, // @[:anonymous source@576.4]
  input          R0_clk, // @[:anonymous source@577.4]
  output [119:0] R0_data, // @[:anonymous source@578.4]
  input          R0_en // @[:anonymous source@579.4]
);
  wire [6:0] mem_0_0_W0_addr; // @[:anonymous source@581.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@581.4]
  wire [29:0] mem_0_0_W0_data; // @[:anonymous source@581.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@581.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@581.4]
  wire [6:0] mem_0_0_R0_addr; // @[:anonymous source@581.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@581.4]
  wire [29:0] mem_0_0_R0_data; // @[:anonymous source@581.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@581.4]
  wire [6:0] mem_0_1_W0_addr; // @[:anonymous source@582.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@582.4]
  wire [29:0] mem_0_1_W0_data; // @[:anonymous source@582.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@582.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@582.4]
  wire [6:0] mem_0_1_R0_addr; // @[:anonymous source@582.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@582.4]
  wire [29:0] mem_0_1_R0_data; // @[:anonymous source@582.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@582.4]
  wire [6:0] mem_0_2_W0_addr; // @[:anonymous source@583.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@583.4]
  wire [29:0] mem_0_2_W0_data; // @[:anonymous source@583.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@583.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@583.4]
  wire [6:0] mem_0_2_R0_addr; // @[:anonymous source@583.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@583.4]
  wire [29:0] mem_0_2_R0_data; // @[:anonymous source@583.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@583.4]
  wire [6:0] mem_0_3_W0_addr; // @[:anonymous source@584.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@584.4]
  wire [29:0] mem_0_3_W0_data; // @[:anonymous source@584.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@584.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@584.4]
  wire [6:0] mem_0_3_R0_addr; // @[:anonymous source@584.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@584.4]
  wire [29:0] mem_0_3_R0_data; // @[:anonymous source@584.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@584.4]
  wire [29:0] R0_data_0_0; // @[:anonymous source@607.4]
  wire [29:0] R0_data_0_1; // @[:anonymous source@611.4]
  wire [29:0] R0_data_0_2; // @[:anonymous source@615.4]
  wire [29:0] R0_data_0_3; // @[:anonymous source@619.4]
  wire [59:0] _GEN_0; // @[:anonymous source@621.4]
  wire [89:0] _GEN_1; // @[:anonymous source@621.4]
  wire [119:0] R0_data_0; // @[:anonymous source@621.4]
  wire [59:0] _GEN_2; // @[:anonymous source@622.4]
  wire [89:0] _GEN_3; // @[:anonymous source@622.4]
  split_meta_0_ext mem_0_0 ( // @[:anonymous source@581.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_meta_0_ext mem_0_1 ( // @[:anonymous source@582.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_meta_0_ext mem_0_2 ( // @[:anonymous source@583.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_meta_0_ext mem_0_3 ( // @[:anonymous source@584.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@607.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@611.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@615.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@619.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@621.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@621.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@621.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@622.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@622.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@622.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@586.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@585.4]
  assign mem_0_0_W0_data = W0_data[29:0]; // @[:anonymous source@587.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@589.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@588.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@606.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@605.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@608.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@591.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@590.4]
  assign mem_0_1_W0_data = W0_data[59:30]; // @[:anonymous source@592.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@594.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@593.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@610.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@609.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@612.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@596.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@595.4]
  assign mem_0_2_W0_data = W0_data[89:60]; // @[:anonymous source@597.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@599.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@598.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@614.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@613.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@616.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@601.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@600.4]
  assign mem_0_3_W0_data = W0_data[119:90]; // @[:anonymous source@602.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@604.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@603.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@618.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@617.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@620.4]
endmodule
module btb_0_ext( // @[:anonymous source@624.2]
  input  [6:0]  W0_addr, // @[:anonymous source@625.4]
  input         W0_clk, // @[:anonymous source@626.4]
  input  [55:0] W0_data, // @[:anonymous source@627.4]
  input         W0_en, // @[:anonymous source@628.4]
  input  [3:0]  W0_mask, // @[:anonymous source@629.4]
  input  [6:0]  R0_addr, // @[:anonymous source@630.4]
  input         R0_clk, // @[:anonymous source@631.4]
  output [55:0] R0_data, // @[:anonymous source@632.4]
  input         R0_en // @[:anonymous source@633.4]
);
  wire [6:0] mem_0_0_W0_addr; // @[:anonymous source@635.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@635.4]
  wire [13:0] mem_0_0_W0_data; // @[:anonymous source@635.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@635.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@635.4]
  wire [6:0] mem_0_0_R0_addr; // @[:anonymous source@635.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@635.4]
  wire [13:0] mem_0_0_R0_data; // @[:anonymous source@635.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@635.4]
  wire [6:0] mem_0_1_W0_addr; // @[:anonymous source@636.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@636.4]
  wire [13:0] mem_0_1_W0_data; // @[:anonymous source@636.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@636.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@636.4]
  wire [6:0] mem_0_1_R0_addr; // @[:anonymous source@636.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@636.4]
  wire [13:0] mem_0_1_R0_data; // @[:anonymous source@636.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@636.4]
  wire [6:0] mem_0_2_W0_addr; // @[:anonymous source@637.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@637.4]
  wire [13:0] mem_0_2_W0_data; // @[:anonymous source@637.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@637.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@637.4]
  wire [6:0] mem_0_2_R0_addr; // @[:anonymous source@637.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@637.4]
  wire [13:0] mem_0_2_R0_data; // @[:anonymous source@637.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@637.4]
  wire [6:0] mem_0_3_W0_addr; // @[:anonymous source@638.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@638.4]
  wire [13:0] mem_0_3_W0_data; // @[:anonymous source@638.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@638.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@638.4]
  wire [6:0] mem_0_3_R0_addr; // @[:anonymous source@638.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@638.4]
  wire [13:0] mem_0_3_R0_data; // @[:anonymous source@638.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@638.4]
  wire [13:0] R0_data_0_0; // @[:anonymous source@661.4]
  wire [13:0] R0_data_0_1; // @[:anonymous source@665.4]
  wire [13:0] R0_data_0_2; // @[:anonymous source@669.4]
  wire [13:0] R0_data_0_3; // @[:anonymous source@673.4]
  wire [27:0] _GEN_0; // @[:anonymous source@675.4]
  wire [41:0] _GEN_1; // @[:anonymous source@675.4]
  wire [55:0] R0_data_0; // @[:anonymous source@675.4]
  wire [27:0] _GEN_2; // @[:anonymous source@676.4]
  wire [41:0] _GEN_3; // @[:anonymous source@676.4]
  split_btb_0_ext mem_0_0 ( // @[:anonymous source@635.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_btb_0_ext mem_0_1 ( // @[:anonymous source@636.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_btb_0_ext mem_0_2 ( // @[:anonymous source@637.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_btb_0_ext mem_0_3 ( // @[:anonymous source@638.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@661.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@665.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@669.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@673.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@675.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@675.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@675.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@676.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@676.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@676.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@640.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@639.4]
  assign mem_0_0_W0_data = W0_data[13:0]; // @[:anonymous source@641.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@643.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@642.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@660.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@659.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@662.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@645.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@644.4]
  assign mem_0_1_W0_data = W0_data[27:14]; // @[:anonymous source@646.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@648.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@647.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@664.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@663.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@666.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@650.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@649.4]
  assign mem_0_2_W0_data = W0_data[41:28]; // @[:anonymous source@651.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@653.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@652.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@668.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@667.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@670.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@655.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@654.4]
  assign mem_0_3_W0_data = W0_data[55:42]; // @[:anonymous source@656.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@658.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@657.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@672.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@671.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@674.4]
endmodule
module ebtb_ext( // @[:anonymous source@678.2]
  input  [6:0]  W0_addr, // @[:anonymous source@679.4]
  input         W0_clk, // @[:anonymous source@680.4]
  input  [39:0] W0_data, // @[:anonymous source@681.4]
  input         W0_en, // @[:anonymous source@682.4]
  input  [6:0]  R0_addr, // @[:anonymous source@683.4]
  input         R0_clk, // @[:anonymous source@684.4]
  output [39:0] R0_data, // @[:anonymous source@685.4]
  input         R0_en // @[:anonymous source@686.4]
);
  wire [6:0] mem_0_0_W0_addr; // @[:anonymous source@688.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@688.4]
  wire [39:0] mem_0_0_W0_data; // @[:anonymous source@688.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@688.4]
  wire [6:0] mem_0_0_R0_addr; // @[:anonymous source@688.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@688.4]
  wire [39:0] mem_0_0_R0_data; // @[:anonymous source@688.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@688.4]
  wire [39:0] R0_data_0_0; // @[:anonymous source@695.4]
  wire [39:0] R0_data_0; // @[:anonymous source@697.4]
  split_ebtb_ext mem_0_0 ( // @[:anonymous source@688.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@695.4]
  assign R0_data_0 = R0_data_0_0; // @[:anonymous source@697.4]
  assign R0_data = mem_0_0_R0_data; // @[:anonymous source@698.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@690.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@689.4]
  assign mem_0_0_W0_data = W0_data; // @[:anonymous source@691.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@692.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@694.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@693.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@696.4]
endmodule
module data_ext( // @[:anonymous source@700.2]
  input  [10:0] W0_addr, // @[:anonymous source@701.4]
  input         W0_clk, // @[:anonymous source@702.4]
  input  [7:0]  W0_data, // @[:anonymous source@703.4]
  input         W0_en, // @[:anonymous source@704.4]
  input  [3:0]  W0_mask, // @[:anonymous source@705.4]
  input  [10:0] R0_addr, // @[:anonymous source@706.4]
  input         R0_clk, // @[:anonymous source@707.4]
  output [7:0]  R0_data, // @[:anonymous source@708.4]
  input         R0_en // @[:anonymous source@709.4]
);
  wire [10:0] mem_0_0_W0_addr; // @[:anonymous source@711.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@711.4]
  wire [1:0] mem_0_0_W0_data; // @[:anonymous source@711.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@711.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@711.4]
  wire [10:0] mem_0_0_R0_addr; // @[:anonymous source@711.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@711.4]
  wire [1:0] mem_0_0_R0_data; // @[:anonymous source@711.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@711.4]
  wire [10:0] mem_0_1_W0_addr; // @[:anonymous source@712.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@712.4]
  wire [1:0] mem_0_1_W0_data; // @[:anonymous source@712.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@712.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@712.4]
  wire [10:0] mem_0_1_R0_addr; // @[:anonymous source@712.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@712.4]
  wire [1:0] mem_0_1_R0_data; // @[:anonymous source@712.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@712.4]
  wire [10:0] mem_0_2_W0_addr; // @[:anonymous source@713.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@713.4]
  wire [1:0] mem_0_2_W0_data; // @[:anonymous source@713.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@713.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@713.4]
  wire [10:0] mem_0_2_R0_addr; // @[:anonymous source@713.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@713.4]
  wire [1:0] mem_0_2_R0_data; // @[:anonymous source@713.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@713.4]
  wire [10:0] mem_0_3_W0_addr; // @[:anonymous source@714.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@714.4]
  wire [1:0] mem_0_3_W0_data; // @[:anonymous source@714.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@714.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@714.4]
  wire [10:0] mem_0_3_R0_addr; // @[:anonymous source@714.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@714.4]
  wire [1:0] mem_0_3_R0_data; // @[:anonymous source@714.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@714.4]
  wire [1:0] R0_data_0_0; // @[:anonymous source@737.4]
  wire [1:0] R0_data_0_1; // @[:anonymous source@741.4]
  wire [1:0] R0_data_0_2; // @[:anonymous source@745.4]
  wire [1:0] R0_data_0_3; // @[:anonymous source@749.4]
  wire [3:0] _GEN_0; // @[:anonymous source@751.4]
  wire [5:0] _GEN_1; // @[:anonymous source@751.4]
  wire [7:0] R0_data_0; // @[:anonymous source@751.4]
  wire [3:0] _GEN_2; // @[:anonymous source@752.4]
  wire [5:0] _GEN_3; // @[:anonymous source@752.4]
  split_data_ext mem_0_0 ( // @[:anonymous source@711.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_data_ext mem_0_1 ( // @[:anonymous source@712.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_data_ext mem_0_2 ( // @[:anonymous source@713.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_data_ext mem_0_3 ( // @[:anonymous source@714.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@737.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@741.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@745.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@749.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@751.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@751.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@751.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@752.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@752.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@752.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@716.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@715.4]
  assign mem_0_0_W0_data = W0_data[1:0]; // @[:anonymous source@717.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@719.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@718.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@736.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@735.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@738.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@721.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@720.4]
  assign mem_0_1_W0_data = W0_data[3:2]; // @[:anonymous source@722.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@724.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@723.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@740.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@739.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@742.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@726.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@725.4]
  assign mem_0_2_W0_data = W0_data[5:4]; // @[:anonymous source@727.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@729.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@728.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@744.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@743.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@746.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@731.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@730.4]
  assign mem_0_3_W0_data = W0_data[7:6]; // @[:anonymous source@732.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@734.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@733.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@748.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@747.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@750.4]
endmodule
module meta_ext( // @[:anonymous source@754.2]
  input  [4:0]   W0_addr, // @[:anonymous source@755.4]
  input          W0_clk, // @[:anonymous source@756.4]
  input  [239:0] W0_data, // @[:anonymous source@757.4]
  input          W0_en, // @[:anonymous source@758.4]
  input  [4:0]   R0_addr, // @[:anonymous source@759.4]
  input          R0_clk, // @[:anonymous source@760.4]
  output [239:0] R0_data, // @[:anonymous source@761.4]
  input          R0_en // @[:anonymous source@762.4]
);
  wire [4:0] mem_0_0_W0_addr; // @[:anonymous source@764.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@764.4]
  wire [239:0] mem_0_0_W0_data; // @[:anonymous source@764.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@764.4]
  wire [4:0] mem_0_0_R0_addr; // @[:anonymous source@764.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@764.4]
  wire [239:0] mem_0_0_R0_data; // @[:anonymous source@764.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@764.4]
  wire [239:0] R0_data_0_0; // @[:anonymous source@771.4]
  wire [239:0] R0_data_0; // @[:anonymous source@773.4]
  split_meta_ext mem_0_0 ( // @[:anonymous source@764.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@771.4]
  assign R0_data_0 = R0_data_0_0; // @[:anonymous source@773.4]
  assign R0_data = mem_0_0_R0_data; // @[:anonymous source@774.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@766.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@765.4]
  assign mem_0_0_W0_data = W0_data; // @[:anonymous source@767.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@768.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@770.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@769.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@772.4]
endmodule
module ghist_0_ext( // @[:anonymous source@776.2]
  input  [4:0]  W0_addr, // @[:anonymous source@777.4]
  input         W0_clk, // @[:anonymous source@778.4]
  input  [71:0] W0_data, // @[:anonymous source@779.4]
  input         W0_en, // @[:anonymous source@780.4]
  input  [4:0]  R0_addr, // @[:anonymous source@781.4]
  input         R0_clk, // @[:anonymous source@782.4]
  output [71:0] R0_data, // @[:anonymous source@783.4]
  input         R0_en // @[:anonymous source@784.4]
);
  wire [4:0] mem_0_0_W0_addr; // @[:anonymous source@786.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@786.4]
  wire [71:0] mem_0_0_W0_data; // @[:anonymous source@786.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@786.4]
  wire [4:0] mem_0_0_R0_addr; // @[:anonymous source@786.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@786.4]
  wire [71:0] mem_0_0_R0_data; // @[:anonymous source@786.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@786.4]
  wire [71:0] R0_data_0_0; // @[:anonymous source@793.4]
  wire [71:0] R0_data_0; // @[:anonymous source@795.4]
  split_ghist_0_ext mem_0_0 ( // @[:anonymous source@786.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@793.4]
  assign R0_data_0 = R0_data_0_0; // @[:anonymous source@795.4]
  assign R0_data = mem_0_0_R0_data; // @[:anonymous source@796.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@788.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@787.4]
  assign mem_0_0_W0_data = W0_data; // @[:anonymous source@789.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@790.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@792.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@791.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@794.4]
endmodule
module rob_debug_inst_mem_ext( // @[:anonymous source@798.2]
  input  [4:0]  W0_addr, // @[:anonymous source@799.4]
  input         W0_clk, // @[:anonymous source@800.4]
  input  [95:0] W0_data, // @[:anonymous source@801.4]
  input         W0_en, // @[:anonymous source@802.4]
  input  [2:0]  W0_mask, // @[:anonymous source@803.4]
  input  [4:0]  R0_addr, // @[:anonymous source@804.4]
  input         R0_clk, // @[:anonymous source@805.4]
  output [95:0] R0_data, // @[:anonymous source@806.4]
  input         R0_en // @[:anonymous source@807.4]
);
  wire [4:0] mem_0_0_W0_addr; // @[:anonymous source@809.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@809.4]
  wire [31:0] mem_0_0_W0_data; // @[:anonymous source@809.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@809.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@809.4]
  wire [4:0] mem_0_0_R0_addr; // @[:anonymous source@809.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@809.4]
  wire [31:0] mem_0_0_R0_data; // @[:anonymous source@809.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@809.4]
  wire [4:0] mem_0_1_W0_addr; // @[:anonymous source@810.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@810.4]
  wire [31:0] mem_0_1_W0_data; // @[:anonymous source@810.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@810.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@810.4]
  wire [4:0] mem_0_1_R0_addr; // @[:anonymous source@810.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@810.4]
  wire [31:0] mem_0_1_R0_data; // @[:anonymous source@810.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@810.4]
  wire [4:0] mem_0_2_W0_addr; // @[:anonymous source@811.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@811.4]
  wire [31:0] mem_0_2_W0_data; // @[:anonymous source@811.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@811.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@811.4]
  wire [4:0] mem_0_2_R0_addr; // @[:anonymous source@811.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@811.4]
  wire [31:0] mem_0_2_R0_data; // @[:anonymous source@811.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@811.4]
  wire [31:0] R0_data_0_0; // @[:anonymous source@829.4]
  wire [31:0] R0_data_0_1; // @[:anonymous source@833.4]
  wire [31:0] R0_data_0_2; // @[:anonymous source@837.4]
  wire [63:0] _GEN_0; // @[:anonymous source@839.4]
  wire [95:0] R0_data_0; // @[:anonymous source@839.4]
  wire [63:0] _GEN_1; // @[:anonymous source@840.4]
  split_rob_debug_inst_mem_ext mem_0_0 ( // @[:anonymous source@809.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_rob_debug_inst_mem_ext mem_0_1 ( // @[:anonymous source@810.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_rob_debug_inst_mem_ext mem_0_2 ( // @[:anonymous source@811.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@829.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@833.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@837.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@839.4]
  assign R0_data_0 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@839.4]
  assign _GEN_1 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@840.4]
  assign R0_data = {R0_data_0_2,_GEN_0}; // @[:anonymous source@840.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@813.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@812.4]
  assign mem_0_0_W0_data = W0_data[31:0]; // @[:anonymous source@814.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@816.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@815.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@828.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@827.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@830.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@818.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@817.4]
  assign mem_0_1_W0_data = W0_data[63:32]; // @[:anonymous source@819.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@821.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@820.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@832.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@831.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@834.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@823.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@822.4]
  assign mem_0_2_W0_data = W0_data[95:64]; // @[:anonymous source@824.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@826.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@825.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@836.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@835.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@838.4]
endmodule
module l2_tlb_ram_ext( // @[:anonymous source@842.2]
  input  [9:0]  RW0_addr, // @[:anonymous source@843.4]
  input         RW0_clk, // @[:anonymous source@844.4]
  input  [43:0] RW0_wdata, // @[:anonymous source@845.4]
  output [43:0] RW0_rdata, // @[:anonymous source@846.4]
  input         RW0_en, // @[:anonymous source@847.4]
  input         RW0_wmode // @[:anonymous source@848.4]
);
  wire [9:0] mem_0_0_RW0_addr; // @[:anonymous source@850.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@850.4]
  wire [43:0] mem_0_0_RW0_wdata; // @[:anonymous source@850.4]
  wire [43:0] mem_0_0_RW0_rdata; // @[:anonymous source@850.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@850.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@850.4]
  wire [43:0] RW0_rdata_0_0; // @[:anonymous source@853.4]
  wire [43:0] RW0_rdata_0; // @[:anonymous source@857.4]
  split_l2_tlb_ram_ext mem_0_0 ( // @[:anonymous source@850.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@853.4]
  assign RW0_rdata_0 = RW0_rdata_0_0; // @[:anonymous source@857.4]
  assign RW0_rdata = mem_0_0_RW0_rdata; // @[:anonymous source@858.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@852.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@851.4]
  assign mem_0_0_RW0_wdata = RW0_wdata; // @[:anonymous source@854.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@856.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@855.4]
endmodule
module split_cc_dir_ext( // @[:anonymous source@860.2]
  input  [9:0]  RW0_addr, // @[:anonymous source@861.4]
  input         RW0_clk, // @[:anonymous source@862.4]
  input  [15:0] RW0_wdata, // @[:anonymous source@863.4]
  output [15:0] RW0_rdata, // @[:anonymous source@864.4]
  input         RW0_en, // @[:anonymous source@865.4]
  input         RW0_wmode, // @[:anonymous source@866.4]
  input         RW0_wmask // @[:anonymous source@867.4]
);
  reg [15:0] ram [0:1023]; // @[:anonymous source@869.4]
  reg [31:0] _RAND_0;
  wire [15:0] ram_RW_0_r_data; // @[:anonymous source@869.4]
  wire [9:0] ram_RW_0_r_addr; // @[:anonymous source@869.4]
  wire [15:0] ram_RW_0_w_data; // @[:anonymous source@869.4]
  wire [9:0] ram_RW_0_w_addr; // @[:anonymous source@869.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@869.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@869.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [9:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@869.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@881.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    ram[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@869.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_cc_banks_0_ext( // @[:anonymous source@884.2]
  input  [12:0] RW0_addr, // @[:anonymous source@885.4]
  input         RW0_clk, // @[:anonymous source@886.4]
  input  [63:0] RW0_wdata, // @[:anonymous source@887.4]
  output [63:0] RW0_rdata, // @[:anonymous source@888.4]
  input         RW0_en, // @[:anonymous source@889.4]
  input         RW0_wmode // @[:anonymous source@890.4]
);
  reg [63:0] ram [0:8191]; // @[:anonymous source@892.4]
  reg [63:0] _RAND_0;
  wire [63:0] ram_RW_0_r_data; // @[:anonymous source@892.4]
  wire [12:0] ram_RW_0_r_addr; // @[:anonymous source@892.4]
  wire [63:0] ram_RW_0_w_data; // @[:anonymous source@892.4]
  wire [12:0] ram_RW_0_w_addr; // @[:anonymous source@892.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@892.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@892.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [12:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@892.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = 1'h1;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@904.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8192; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[12:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@892.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_tag_array_ext( // @[:anonymous source@907.2]
  input  [5:0]  RW0_addr, // @[:anonymous source@908.4]
  input         RW0_clk, // @[:anonymous source@909.4]
  input  [21:0] RW0_wdata, // @[:anonymous source@910.4]
  output [21:0] RW0_rdata, // @[:anonymous source@911.4]
  input         RW0_en, // @[:anonymous source@912.4]
  input         RW0_wmode, // @[:anonymous source@913.4]
  input         RW0_wmask // @[:anonymous source@914.4]
);
  reg [21:0] ram [0:63]; // @[:anonymous source@916.4]
  reg [31:0] _RAND_0;
  wire [21:0] ram_RW_0_r_data; // @[:anonymous source@916.4]
  wire [5:0] ram_RW_0_r_addr; // @[:anonymous source@916.4]
  wire [21:0] ram_RW_0_w_data; // @[:anonymous source@916.4]
  wire [5:0] ram_RW_0_w_addr; // @[:anonymous source@916.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@916.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@916.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [5:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@916.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@928.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram[initvar] = _RAND_0[21:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@916.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_array_0_0_ext( // @[:anonymous source@931.2]
  input  [7:0]  W0_addr, // @[:anonymous source@932.4]
  input         W0_clk, // @[:anonymous source@933.4]
  input  [63:0] W0_data, // @[:anonymous source@934.4]
  input         W0_en, // @[:anonymous source@935.4]
  input         W0_mask, // @[:anonymous source@936.4]
  input  [7:0]  R0_addr, // @[:anonymous source@937.4]
  input         R0_clk, // @[:anonymous source@938.4]
  output [63:0] R0_data, // @[:anonymous source@939.4]
  input         R0_en // @[:anonymous source@940.4]
);
  reg [63:0] ram [0:255]; // @[:anonymous source@942.4]
  reg [63:0] _RAND_0;
  wire [63:0] ram_R_0_data; // @[:anonymous source@942.4]
  wire [7:0] ram_R_0_addr; // @[:anonymous source@942.4]
  wire [63:0] ram_W_0_data; // @[:anonymous source@942.4]
  wire [7:0] ram_W_0_addr; // @[:anonymous source@942.4]
  wire  ram_W_0_mask; // @[:anonymous source@942.4]
  wire  ram_W_0_en; // @[:anonymous source@942.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [7:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@942.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@953.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@942.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_tag_array_0_ext( // @[:anonymous source@960.2]
  input  [5:0]  RW0_addr, // @[:anonymous source@961.4]
  input         RW0_clk, // @[:anonymous source@962.4]
  input  [19:0] RW0_wdata, // @[:anonymous source@963.4]
  output [19:0] RW0_rdata, // @[:anonymous source@964.4]
  input         RW0_en, // @[:anonymous source@965.4]
  input         RW0_wmode, // @[:anonymous source@966.4]
  input         RW0_wmask // @[:anonymous source@967.4]
);
  reg [19:0] ram [0:63]; // @[:anonymous source@969.4]
  reg [31:0] _RAND_0;
  wire [19:0] ram_RW_0_r_data; // @[:anonymous source@969.4]
  wire [5:0] ram_RW_0_r_addr; // @[:anonymous source@969.4]
  wire [19:0] ram_RW_0_w_data; // @[:anonymous source@969.4]
  wire [5:0] ram_RW_0_w_addr; // @[:anonymous source@969.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@969.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@969.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [5:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@969.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@981.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram[initvar] = _RAND_0[19:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@969.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_dataArrayB0Way_0_ext( // @[:anonymous source@984.2]
  input  [7:0]  RW0_addr, // @[:anonymous source@985.4]
  input         RW0_clk, // @[:anonymous source@986.4]
  input  [63:0] RW0_wdata, // @[:anonymous source@987.4]
  output [63:0] RW0_rdata, // @[:anonymous source@988.4]
  input         RW0_en, // @[:anonymous source@989.4]
  input         RW0_wmode // @[:anonymous source@990.4]
);
  reg [63:0] ram [0:255]; // @[:anonymous source@992.4]
  reg [63:0] _RAND_0;
  wire [63:0] ram_RW_0_r_data; // @[:anonymous source@992.4]
  wire [7:0] ram_RW_0_r_addr; // @[:anonymous source@992.4]
  wire [63:0] ram_RW_0_w_data; // @[:anonymous source@992.4]
  wire [7:0] ram_RW_0_w_addr; // @[:anonymous source@992.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@992.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@992.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [7:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@992.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = 1'h1;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@1004.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@992.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_hi_us_ext( // @[:anonymous source@1007.2]
  input  [6:0] W0_addr, // @[:anonymous source@1008.4]
  input        W0_clk, // @[:anonymous source@1009.4]
  input        W0_data, // @[:anonymous source@1010.4]
  input        W0_en, // @[:anonymous source@1011.4]
  input        W0_mask, // @[:anonymous source@1012.4]
  input  [6:0] R0_addr, // @[:anonymous source@1013.4]
  input        R0_clk, // @[:anonymous source@1014.4]
  output       R0_data, // @[:anonymous source@1015.4]
  input        R0_en // @[:anonymous source@1016.4]
);
  reg  ram [0:127]; // @[:anonymous source@1018.4]
  reg [31:0] _RAND_0;
  wire  ram_R_0_data; // @[:anonymous source@1018.4]
  wire [6:0] ram_R_0_addr; // @[:anonymous source@1018.4]
  wire  ram_W_0_data; // @[:anonymous source@1018.4]
  wire [6:0] ram_W_0_addr; // @[:anonymous source@1018.4]
  wire  ram_W_0_mask; // @[:anonymous source@1018.4]
  wire  ram_W_0_en; // @[:anonymous source@1018.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1018.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1029.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1018.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_table_ext( // @[:anonymous source@1036.2]
  input  [6:0]  W0_addr, // @[:anonymous source@1037.4]
  input         W0_clk, // @[:anonymous source@1038.4]
  input  [10:0] W0_data, // @[:anonymous source@1039.4]
  input         W0_en, // @[:anonymous source@1040.4]
  input         W0_mask, // @[:anonymous source@1041.4]
  input  [6:0]  R0_addr, // @[:anonymous source@1042.4]
  input         R0_clk, // @[:anonymous source@1043.4]
  output [10:0] R0_data, // @[:anonymous source@1044.4]
  input         R0_en // @[:anonymous source@1045.4]
);
  reg [10:0] ram [0:127]; // @[:anonymous source@1047.4]
  reg [31:0] _RAND_0;
  wire [10:0] ram_R_0_data; // @[:anonymous source@1047.4]
  wire [6:0] ram_R_0_addr; // @[:anonymous source@1047.4]
  wire [10:0] ram_W_0_data; // @[:anonymous source@1047.4]
  wire [6:0] ram_W_0_addr; // @[:anonymous source@1047.4]
  wire  ram_W_0_mask; // @[:anonymous source@1047.4]
  wire  ram_W_0_en; // @[:anonymous source@1047.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1047.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1058.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[10:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1047.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_hi_us_0_ext( // @[:anonymous source@1065.2]
  input  [7:0] W0_addr, // @[:anonymous source@1066.4]
  input        W0_clk, // @[:anonymous source@1067.4]
  input        W0_data, // @[:anonymous source@1068.4]
  input        W0_en, // @[:anonymous source@1069.4]
  input        W0_mask, // @[:anonymous source@1070.4]
  input  [7:0] R0_addr, // @[:anonymous source@1071.4]
  input        R0_clk, // @[:anonymous source@1072.4]
  output       R0_data, // @[:anonymous source@1073.4]
  input        R0_en // @[:anonymous source@1074.4]
);
  reg  ram [0:255]; // @[:anonymous source@1076.4]
  reg [31:0] _RAND_0;
  wire  ram_R_0_data; // @[:anonymous source@1076.4]
  wire [7:0] ram_R_0_addr; // @[:anonymous source@1076.4]
  wire  ram_W_0_data; // @[:anonymous source@1076.4]
  wire [7:0] ram_W_0_addr; // @[:anonymous source@1076.4]
  wire  ram_W_0_mask; // @[:anonymous source@1076.4]
  wire  ram_W_0_en; // @[:anonymous source@1076.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [7:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1076.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1087.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1076.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_table_0_ext( // @[:anonymous source@1094.2]
  input  [7:0]  W0_addr, // @[:anonymous source@1095.4]
  input         W0_clk, // @[:anonymous source@1096.4]
  input  [11:0] W0_data, // @[:anonymous source@1097.4]
  input         W0_en, // @[:anonymous source@1098.4]
  input         W0_mask, // @[:anonymous source@1099.4]
  input  [7:0]  R0_addr, // @[:anonymous source@1100.4]
  input         R0_clk, // @[:anonymous source@1101.4]
  output [11:0] R0_data, // @[:anonymous source@1102.4]
  input         R0_en // @[:anonymous source@1103.4]
);
  reg [11:0] ram [0:255]; // @[:anonymous source@1105.4]
  reg [31:0] _RAND_0;
  wire [11:0] ram_R_0_data; // @[:anonymous source@1105.4]
  wire [7:0] ram_R_0_addr; // @[:anonymous source@1105.4]
  wire [11:0] ram_W_0_data; // @[:anonymous source@1105.4]
  wire [7:0] ram_W_0_addr; // @[:anonymous source@1105.4]
  wire  ram_W_0_mask; // @[:anonymous source@1105.4]
  wire  ram_W_0_en; // @[:anonymous source@1105.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [7:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1105.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1116.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram[initvar] = _RAND_0[11:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1105.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_table_1_ext( // @[:anonymous source@1123.2]
  input  [6:0]  W0_addr, // @[:anonymous source@1124.4]
  input         W0_clk, // @[:anonymous source@1125.4]
  input  [12:0] W0_data, // @[:anonymous source@1126.4]
  input         W0_en, // @[:anonymous source@1127.4]
  input         W0_mask, // @[:anonymous source@1128.4]
  input  [6:0]  R0_addr, // @[:anonymous source@1129.4]
  input         R0_clk, // @[:anonymous source@1130.4]
  output [12:0] R0_data, // @[:anonymous source@1131.4]
  input         R0_en // @[:anonymous source@1132.4]
);
  reg [12:0] ram [0:127]; // @[:anonymous source@1134.4]
  reg [31:0] _RAND_0;
  wire [12:0] ram_R_0_data; // @[:anonymous source@1134.4]
  wire [6:0] ram_R_0_addr; // @[:anonymous source@1134.4]
  wire [12:0] ram_W_0_data; // @[:anonymous source@1134.4]
  wire [6:0] ram_W_0_addr; // @[:anonymous source@1134.4]
  wire  ram_W_0_mask; // @[:anonymous source@1134.4]
  wire  ram_W_0_en; // @[:anonymous source@1134.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1134.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1145.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[12:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1134.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_meta_0_ext( // @[:anonymous source@1152.2]
  input  [6:0]  W0_addr, // @[:anonymous source@1153.4]
  input         W0_clk, // @[:anonymous source@1154.4]
  input  [29:0] W0_data, // @[:anonymous source@1155.4]
  input         W0_en, // @[:anonymous source@1156.4]
  input         W0_mask, // @[:anonymous source@1157.4]
  input  [6:0]  R0_addr, // @[:anonymous source@1158.4]
  input         R0_clk, // @[:anonymous source@1159.4]
  output [29:0] R0_data, // @[:anonymous source@1160.4]
  input         R0_en // @[:anonymous source@1161.4]
);
  reg [29:0] ram [0:127]; // @[:anonymous source@1163.4]
  reg [31:0] _RAND_0;
  wire [29:0] ram_R_0_data; // @[:anonymous source@1163.4]
  wire [6:0] ram_R_0_addr; // @[:anonymous source@1163.4]
  wire [29:0] ram_W_0_data; // @[:anonymous source@1163.4]
  wire [6:0] ram_W_0_addr; // @[:anonymous source@1163.4]
  wire  ram_W_0_mask; // @[:anonymous source@1163.4]
  wire  ram_W_0_en; // @[:anonymous source@1163.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1163.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1174.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[29:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1163.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_btb_0_ext( // @[:anonymous source@1181.2]
  input  [6:0]  W0_addr, // @[:anonymous source@1182.4]
  input         W0_clk, // @[:anonymous source@1183.4]
  input  [13:0] W0_data, // @[:anonymous source@1184.4]
  input         W0_en, // @[:anonymous source@1185.4]
  input         W0_mask, // @[:anonymous source@1186.4]
  input  [6:0]  R0_addr, // @[:anonymous source@1187.4]
  input         R0_clk, // @[:anonymous source@1188.4]
  output [13:0] R0_data, // @[:anonymous source@1189.4]
  input         R0_en // @[:anonymous source@1190.4]
);
  reg [13:0] ram [0:127]; // @[:anonymous source@1192.4]
  reg [31:0] _RAND_0;
  wire [13:0] ram_R_0_data; // @[:anonymous source@1192.4]
  wire [6:0] ram_R_0_addr; // @[:anonymous source@1192.4]
  wire [13:0] ram_W_0_data; // @[:anonymous source@1192.4]
  wire [6:0] ram_W_0_addr; // @[:anonymous source@1192.4]
  wire  ram_W_0_mask; // @[:anonymous source@1192.4]
  wire  ram_W_0_en; // @[:anonymous source@1192.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1192.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1203.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[13:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1192.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_ebtb_ext( // @[:anonymous source@1210.2]
  input  [6:0]  W0_addr, // @[:anonymous source@1211.4]
  input         W0_clk, // @[:anonymous source@1212.4]
  input  [39:0] W0_data, // @[:anonymous source@1213.4]
  input         W0_en, // @[:anonymous source@1214.4]
  input  [6:0]  R0_addr, // @[:anonymous source@1215.4]
  input         R0_clk, // @[:anonymous source@1216.4]
  output [39:0] R0_data, // @[:anonymous source@1217.4]
  input         R0_en // @[:anonymous source@1218.4]
);
  reg [39:0] ram [0:127]; // @[:anonymous source@1220.4]
  reg [63:0] _RAND_0;
  wire [39:0] ram_R_0_data; // @[:anonymous source@1220.4]
  wire [6:0] ram_R_0_addr; // @[:anonymous source@1220.4]
  wire [39:0] ram_W_0_data; // @[:anonymous source@1220.4]
  wire [6:0] ram_W_0_addr; // @[:anonymous source@1220.4]
  wire  ram_W_0_mask; // @[:anonymous source@1220.4]
  wire  ram_W_0_en; // @[:anonymous source@1220.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1220.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = 1'h1;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1231.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[39:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1220.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_data_ext( // @[:anonymous source@1238.2]
  input  [10:0] W0_addr, // @[:anonymous source@1239.4]
  input         W0_clk, // @[:anonymous source@1240.4]
  input  [1:0]  W0_data, // @[:anonymous source@1241.4]
  input         W0_en, // @[:anonymous source@1242.4]
  input         W0_mask, // @[:anonymous source@1243.4]
  input  [10:0] R0_addr, // @[:anonymous source@1244.4]
  input         R0_clk, // @[:anonymous source@1245.4]
  output [1:0]  R0_data, // @[:anonymous source@1246.4]
  input         R0_en // @[:anonymous source@1247.4]
);
  reg [1:0] ram [0:2047]; // @[:anonymous source@1249.4]
  reg [31:0] _RAND_0;
  wire [1:0] ram_R_0_data; // @[:anonymous source@1249.4]
  wire [10:0] ram_R_0_addr; // @[:anonymous source@1249.4]
  wire [1:0] ram_W_0_data; // @[:anonymous source@1249.4]
  wire [10:0] ram_W_0_addr; // @[:anonymous source@1249.4]
  wire  ram_W_0_mask; // @[:anonymous source@1249.4]
  wire  ram_W_0_en; // @[:anonymous source@1249.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [10:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1249.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1260.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    ram[initvar] = _RAND_0[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[10:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1249.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_meta_ext( // @[:anonymous source@1267.2]
  input  [4:0]   W0_addr, // @[:anonymous source@1268.4]
  input          W0_clk, // @[:anonymous source@1269.4]
  input  [239:0] W0_data, // @[:anonymous source@1270.4]
  input          W0_en, // @[:anonymous source@1271.4]
  input  [4:0]   R0_addr, // @[:anonymous source@1272.4]
  input          R0_clk, // @[:anonymous source@1273.4]
  output [239:0] R0_data, // @[:anonymous source@1274.4]
  input          R0_en // @[:anonymous source@1275.4]
);
  reg [239:0] ram [0:31]; // @[:anonymous source@1277.4]
  reg [255:0] _RAND_0;
  wire [239:0] ram_R_0_data; // @[:anonymous source@1277.4]
  wire [4:0] ram_R_0_addr; // @[:anonymous source@1277.4]
  wire [239:0] ram_W_0_data; // @[:anonymous source@1277.4]
  wire [4:0] ram_W_0_addr; // @[:anonymous source@1277.4]
  wire  ram_W_0_mask; // @[:anonymous source@1277.4]
  wire  ram_W_0_en; // @[:anonymous source@1277.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [4:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1277.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = 1'h1;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1288.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {8{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    ram[initvar] = _RAND_0[239:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1277.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_ghist_0_ext( // @[:anonymous source@1295.2]
  input  [4:0]  W0_addr, // @[:anonymous source@1296.4]
  input         W0_clk, // @[:anonymous source@1297.4]
  input  [71:0] W0_data, // @[:anonymous source@1298.4]
  input         W0_en, // @[:anonymous source@1299.4]
  input  [4:0]  R0_addr, // @[:anonymous source@1300.4]
  input         R0_clk, // @[:anonymous source@1301.4]
  output [71:0] R0_data, // @[:anonymous source@1302.4]
  input         R0_en // @[:anonymous source@1303.4]
);
  reg [71:0] ram [0:31]; // @[:anonymous source@1305.4]
  reg [95:0] _RAND_0;
  wire [71:0] ram_R_0_data; // @[:anonymous source@1305.4]
  wire [4:0] ram_R_0_addr; // @[:anonymous source@1305.4]
  wire [71:0] ram_W_0_data; // @[:anonymous source@1305.4]
  wire [4:0] ram_W_0_addr; // @[:anonymous source@1305.4]
  wire  ram_W_0_mask; // @[:anonymous source@1305.4]
  wire  ram_W_0_en; // @[:anonymous source@1305.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [4:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1305.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = 1'h1;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1316.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {3{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    ram[initvar] = _RAND_0[71:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1305.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_rob_debug_inst_mem_ext( // @[:anonymous source@1323.2]
  input  [4:0]  W0_addr, // @[:anonymous source@1324.4]
  input         W0_clk, // @[:anonymous source@1325.4]
  input  [31:0] W0_data, // @[:anonymous source@1326.4]
  input         W0_en, // @[:anonymous source@1327.4]
  input         W0_mask, // @[:anonymous source@1328.4]
  input  [4:0]  R0_addr, // @[:anonymous source@1329.4]
  input         R0_clk, // @[:anonymous source@1330.4]
  output [31:0] R0_data, // @[:anonymous source@1331.4]
  input         R0_en // @[:anonymous source@1332.4]
);
  reg [31:0] ram [0:31]; // @[:anonymous source@1334.4]
  reg [31:0] _RAND_0;
  wire [31:0] ram_R_0_data; // @[:anonymous source@1334.4]
  wire [4:0] ram_R_0_addr; // @[:anonymous source@1334.4]
  wire [31:0] ram_W_0_data; // @[:anonymous source@1334.4]
  wire [4:0] ram_W_0_addr; // @[:anonymous source@1334.4]
  wire  ram_W_0_mask; // @[:anonymous source@1334.4]
  wire  ram_W_0_en; // @[:anonymous source@1334.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [4:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1334.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1345.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    ram[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1334.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_l2_tlb_ram_ext( // @[:anonymous source@1352.2]
  input  [9:0]  RW0_addr, // @[:anonymous source@1353.4]
  input         RW0_clk, // @[:anonymous source@1354.4]
  input  [43:0] RW0_wdata, // @[:anonymous source@1355.4]
  output [43:0] RW0_rdata, // @[:anonymous source@1356.4]
  input         RW0_en, // @[:anonymous source@1357.4]
  input         RW0_wmode // @[:anonymous source@1358.4]
);
  reg [43:0] ram [0:1023]; // @[:anonymous source@1360.4]
  reg [63:0] _RAND_0;
  wire [43:0] ram_RW_0_r_data; // @[:anonymous source@1360.4]
  wire [9:0] ram_RW_0_r_addr; // @[:anonymous source@1360.4]
  wire [43:0] ram_RW_0_w_data; // @[:anonymous source@1360.4]
  wire [9:0] ram_RW_0_w_addr; // @[:anonymous source@1360.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@1360.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@1360.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [9:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@1360.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = 1'h1;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@1372.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    ram[initvar] = _RAND_0[43:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@1360.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
